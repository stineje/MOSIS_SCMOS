library IEEE; 
use IEEE.std_logic_1164.all;

entity Dadda53 is
	port(	Y : in  std_logic_vector(51 downto 0);
		X : in  std_logic_vector(51 downto 0);
		S : out std_logic_vector(105 downto 0);
		C : out std_logic_vector(105 downto 0));
end Dadda53;

architecture Structure of Dadda53 is

component and2
	port(	X : in  std_logic;
		Y : in  std_logic;
		O : out std_logic);
end component;

component full_adder 
	port(	A : in  std_logic;
                B : in  std_logic;
		CIN : in  std_logic;
		S : out std_logic;
                COUT : out std_logic);
end component;

component half_adder 
	port(	A : in  std_logic;
		CIN : in  std_logic;
		S : out std_logic;
                COUT : out std_logic);
end component;

	signal N0_0_0 : std_logic;
	signal N0_0_1 : std_logic;
	signal N0_0_2 : std_logic;
	signal N0_0_3 : std_logic;
	signal N0_0_4 : std_logic;
	signal N0_0_5 : std_logic;
	signal N0_0_6 : std_logic;
	signal N0_0_7 : std_logic;
	signal N0_0_8 : std_logic;
	signal N0_0_9 : std_logic;
	signal N0_0_10 : std_logic;
	signal N0_0_11 : std_logic;
	signal N0_0_12 : std_logic;
	signal N0_0_13 : std_logic;
	signal N0_0_14 : std_logic;
	signal N0_0_15 : std_logic;
	signal N0_0_16 : std_logic;
	signal N0_0_17 : std_logic;
	signal N0_0_18 : std_logic;
	signal N0_0_19 : std_logic;
	signal N0_0_20 : std_logic;
	signal N0_0_21 : std_logic;
	signal N0_0_22 : std_logic;
	signal N0_0_23 : std_logic;
	signal N0_0_24 : std_logic;
	signal N0_0_25 : std_logic;
	signal N0_0_26 : std_logic;
	signal N0_0_27 : std_logic;
	signal N0_0_28 : std_logic;
	signal N0_0_29 : std_logic;
	signal N0_0_30 : std_logic;
	signal N0_0_31 : std_logic;
	signal N0_0_32 : std_logic;
	signal N0_0_33 : std_logic;
	signal N0_0_34 : std_logic;
	signal N0_0_35 : std_logic;
	signal N0_0_36 : std_logic;
	signal N0_0_37 : std_logic;
	signal N0_0_38 : std_logic;
	signal N0_0_39 : std_logic;
	signal N0_0_40 : std_logic;
	signal N0_0_41 : std_logic;
	signal N0_0_42 : std_logic;
	signal N0_0_43 : std_logic;
	signal N0_0_44 : std_logic;
	signal N0_0_45 : std_logic;
	signal N0_0_46 : std_logic;
	signal N0_0_47 : std_logic;
	signal N0_0_48 : std_logic;
	signal N0_0_49 : std_logic;
	signal N0_0_50 : std_logic;
	signal N0_0_51 : std_logic;
	signal N0_0_52 : std_logic;
	signal N0_1_1 : std_logic;
	signal N0_1_2 : std_logic;
	signal N0_1_3 : std_logic;
	signal N0_1_4 : std_logic;
	signal N0_1_5 : std_logic;
	signal N0_1_6 : std_logic;
	signal N0_1_7 : std_logic;
	signal N0_1_8 : std_logic;
	signal N0_1_9 : std_logic;
	signal N0_1_10 : std_logic;
	signal N0_1_11 : std_logic;
	signal N0_1_12 : std_logic;
	signal N0_1_13 : std_logic;
	signal N0_1_14 : std_logic;
	signal N0_1_15 : std_logic;
	signal N0_1_16 : std_logic;
	signal N0_1_17 : std_logic;
	signal N0_1_18 : std_logic;
	signal N0_1_19 : std_logic;
	signal N0_1_20 : std_logic;
	signal N0_1_21 : std_logic;
	signal N0_1_22 : std_logic;
	signal N0_1_23 : std_logic;
	signal N0_1_24 : std_logic;
	signal N0_1_25 : std_logic;
	signal N0_1_26 : std_logic;
	signal N0_1_27 : std_logic;
	signal N0_1_28 : std_logic;
	signal N0_1_29 : std_logic;
	signal N0_1_30 : std_logic;
	signal N0_1_31 : std_logic;
	signal N0_1_32 : std_logic;
	signal N0_1_33 : std_logic;
	signal N0_1_34 : std_logic;
	signal N0_1_35 : std_logic;
	signal N0_1_36 : std_logic;
	signal N0_1_37 : std_logic;
	signal N0_1_38 : std_logic;
	signal N0_1_39 : std_logic;
	signal N0_1_40 : std_logic;
	signal N0_1_41 : std_logic;
	signal N0_1_42 : std_logic;
	signal N0_1_43 : std_logic;
	signal N0_1_44 : std_logic;
	signal N0_1_45 : std_logic;
	signal N0_1_46 : std_logic;
	signal N0_1_47 : std_logic;
	signal N0_1_48 : std_logic;
	signal N0_1_49 : std_logic;
	signal N0_1_50 : std_logic;
	signal N0_1_51 : std_logic;
	signal N0_1_52 : std_logic;
	signal N0_1_53 : std_logic;
	signal N0_2_2 : std_logic;
	signal N0_2_3 : std_logic;
	signal N0_2_4 : std_logic;
	signal N0_2_5 : std_logic;
	signal N0_2_6 : std_logic;
	signal N0_2_7 : std_logic;
	signal N0_2_8 : std_logic;
	signal N0_2_9 : std_logic;
	signal N0_2_10 : std_logic;
	signal N0_2_11 : std_logic;
	signal N0_2_12 : std_logic;
	signal N0_2_13 : std_logic;
	signal N0_2_14 : std_logic;
	signal N0_2_15 : std_logic;
	signal N0_2_16 : std_logic;
	signal N0_2_17 : std_logic;
	signal N0_2_18 : std_logic;
	signal N0_2_19 : std_logic;
	signal N0_2_20 : std_logic;
	signal N0_2_21 : std_logic;
	signal N0_2_22 : std_logic;
	signal N0_2_23 : std_logic;
	signal N0_2_24 : std_logic;
	signal N0_2_25 : std_logic;
	signal N0_2_26 : std_logic;
	signal N0_2_27 : std_logic;
	signal N0_2_28 : std_logic;
	signal N0_2_29 : std_logic;
	signal N0_2_30 : std_logic;
	signal N0_2_31 : std_logic;
	signal N0_2_32 : std_logic;
	signal N0_2_33 : std_logic;
	signal N0_2_34 : std_logic;
	signal N0_2_35 : std_logic;
	signal N0_2_36 : std_logic;
	signal N0_2_37 : std_logic;
	signal N0_2_38 : std_logic;
	signal N0_2_39 : std_logic;
	signal N0_2_40 : std_logic;
	signal N0_2_41 : std_logic;
	signal N0_2_42 : std_logic;
	signal N0_2_43 : std_logic;
	signal N0_2_44 : std_logic;
	signal N0_2_45 : std_logic;
	signal N0_2_46 : std_logic;
	signal N0_2_47 : std_logic;
	signal N0_2_48 : std_logic;
	signal N0_2_49 : std_logic;
	signal N0_2_50 : std_logic;
	signal N0_2_51 : std_logic;
	signal N0_2_52 : std_logic;
	signal N0_2_53 : std_logic;
	signal N0_2_54 : std_logic;
	signal N0_3_3 : std_logic;
	signal N0_3_4 : std_logic;
	signal N0_3_5 : std_logic;
	signal N0_3_6 : std_logic;
	signal N0_3_7 : std_logic;
	signal N0_3_8 : std_logic;
	signal N0_3_9 : std_logic;
	signal N0_3_10 : std_logic;
	signal N0_3_11 : std_logic;
	signal N0_3_12 : std_logic;
	signal N0_3_13 : std_logic;
	signal N0_3_14 : std_logic;
	signal N0_3_15 : std_logic;
	signal N0_3_16 : std_logic;
	signal N0_3_17 : std_logic;
	signal N0_3_18 : std_logic;
	signal N0_3_19 : std_logic;
	signal N0_3_20 : std_logic;
	signal N0_3_21 : std_logic;
	signal N0_3_22 : std_logic;
	signal N0_3_23 : std_logic;
	signal N0_3_24 : std_logic;
	signal N0_3_25 : std_logic;
	signal N0_3_26 : std_logic;
	signal N0_3_27 : std_logic;
	signal N0_3_28 : std_logic;
	signal N0_3_29 : std_logic;
	signal N0_3_30 : std_logic;
	signal N0_3_31 : std_logic;
	signal N0_3_32 : std_logic;
	signal N0_3_33 : std_logic;
	signal N0_3_34 : std_logic;
	signal N0_3_35 : std_logic;
	signal N0_3_36 : std_logic;
	signal N0_3_37 : std_logic;
	signal N0_3_38 : std_logic;
	signal N0_3_39 : std_logic;
	signal N0_3_40 : std_logic;
	signal N0_3_41 : std_logic;
	signal N0_3_42 : std_logic;
	signal N0_3_43 : std_logic;
	signal N0_3_44 : std_logic;
	signal N0_3_45 : std_logic;
	signal N0_3_46 : std_logic;
	signal N0_3_47 : std_logic;
	signal N0_3_48 : std_logic;
	signal N0_3_49 : std_logic;
	signal N0_3_50 : std_logic;
	signal N0_3_51 : std_logic;
	signal N0_3_52 : std_logic;
	signal N0_3_53 : std_logic;
	signal N0_3_54 : std_logic;
	signal N0_3_55 : std_logic;
	signal N0_4_4 : std_logic;
	signal N0_4_5 : std_logic;
	signal N0_4_6 : std_logic;
	signal N0_4_7 : std_logic;
	signal N0_4_8 : std_logic;
	signal N0_4_9 : std_logic;
	signal N0_4_10 : std_logic;
	signal N0_4_11 : std_logic;
	signal N0_4_12 : std_logic;
	signal N0_4_13 : std_logic;
	signal N0_4_14 : std_logic;
	signal N0_4_15 : std_logic;
	signal N0_4_16 : std_logic;
	signal N0_4_17 : std_logic;
	signal N0_4_18 : std_logic;
	signal N0_4_19 : std_logic;
	signal N0_4_20 : std_logic;
	signal N0_4_21 : std_logic;
	signal N0_4_22 : std_logic;
	signal N0_4_23 : std_logic;
	signal N0_4_24 : std_logic;
	signal N0_4_25 : std_logic;
	signal N0_4_26 : std_logic;
	signal N0_4_27 : std_logic;
	signal N0_4_28 : std_logic;
	signal N0_4_29 : std_logic;
	signal N0_4_30 : std_logic;
	signal N0_4_31 : std_logic;
	signal N0_4_32 : std_logic;
	signal N0_4_33 : std_logic;
	signal N0_4_34 : std_logic;
	signal N0_4_35 : std_logic;
	signal N0_4_36 : std_logic;
	signal N0_4_37 : std_logic;
	signal N0_4_38 : std_logic;
	signal N0_4_39 : std_logic;
	signal N0_4_40 : std_logic;
	signal N0_4_41 : std_logic;
	signal N0_4_42 : std_logic;
	signal N0_4_43 : std_logic;
	signal N0_4_44 : std_logic;
	signal N0_4_45 : std_logic;
	signal N0_4_46 : std_logic;
	signal N0_4_47 : std_logic;
	signal N0_4_48 : std_logic;
	signal N0_4_49 : std_logic;
	signal N0_4_50 : std_logic;
	signal N0_4_51 : std_logic;
	signal N0_4_52 : std_logic;
	signal N0_4_53 : std_logic;
	signal N0_4_54 : std_logic;
	signal N0_4_55 : std_logic;
	signal N0_4_56 : std_logic;
	signal N0_5_5 : std_logic;
	signal N0_5_6 : std_logic;
	signal N0_5_7 : std_logic;
	signal N0_5_8 : std_logic;
	signal N0_5_9 : std_logic;
	signal N0_5_10 : std_logic;
	signal N0_5_11 : std_logic;
	signal N0_5_12 : std_logic;
	signal N0_5_13 : std_logic;
	signal N0_5_14 : std_logic;
	signal N0_5_15 : std_logic;
	signal N0_5_16 : std_logic;
	signal N0_5_17 : std_logic;
	signal N0_5_18 : std_logic;
	signal N0_5_19 : std_logic;
	signal N0_5_20 : std_logic;
	signal N0_5_21 : std_logic;
	signal N0_5_22 : std_logic;
	signal N0_5_23 : std_logic;
	signal N0_5_24 : std_logic;
	signal N0_5_25 : std_logic;
	signal N0_5_26 : std_logic;
	signal N0_5_27 : std_logic;
	signal N0_5_28 : std_logic;
	signal N0_5_29 : std_logic;
	signal N0_5_30 : std_logic;
	signal N0_5_31 : std_logic;
	signal N0_5_32 : std_logic;
	signal N0_5_33 : std_logic;
	signal N0_5_34 : std_logic;
	signal N0_5_35 : std_logic;
	signal N0_5_36 : std_logic;
	signal N0_5_37 : std_logic;
	signal N0_5_38 : std_logic;
	signal N0_5_39 : std_logic;
	signal N0_5_40 : std_logic;
	signal N0_5_41 : std_logic;
	signal N0_5_42 : std_logic;
	signal N0_5_43 : std_logic;
	signal N0_5_44 : std_logic;
	signal N0_5_45 : std_logic;
	signal N0_5_46 : std_logic;
	signal N0_5_47 : std_logic;
	signal N0_5_48 : std_logic;
	signal N0_5_49 : std_logic;
	signal N0_5_50 : std_logic;
	signal N0_5_51 : std_logic;
	signal N0_5_52 : std_logic;
	signal N0_5_53 : std_logic;
	signal N0_5_54 : std_logic;
	signal N0_5_55 : std_logic;
	signal N0_5_56 : std_logic;
	signal N0_5_57 : std_logic;
	signal N0_6_6 : std_logic;
	signal N0_6_7 : std_logic;
	signal N0_6_8 : std_logic;
	signal N0_6_9 : std_logic;
	signal N0_6_10 : std_logic;
	signal N0_6_11 : std_logic;
	signal N0_6_12 : std_logic;
	signal N0_6_13 : std_logic;
	signal N0_6_14 : std_logic;
	signal N0_6_15 : std_logic;
	signal N0_6_16 : std_logic;
	signal N0_6_17 : std_logic;
	signal N0_6_18 : std_logic;
	signal N0_6_19 : std_logic;
	signal N0_6_20 : std_logic;
	signal N0_6_21 : std_logic;
	signal N0_6_22 : std_logic;
	signal N0_6_23 : std_logic;
	signal N0_6_24 : std_logic;
	signal N0_6_25 : std_logic;
	signal N0_6_26 : std_logic;
	signal N0_6_27 : std_logic;
	signal N0_6_28 : std_logic;
	signal N0_6_29 : std_logic;
	signal N0_6_30 : std_logic;
	signal N0_6_31 : std_logic;
	signal N0_6_32 : std_logic;
	signal N0_6_33 : std_logic;
	signal N0_6_34 : std_logic;
	signal N0_6_35 : std_logic;
	signal N0_6_36 : std_logic;
	signal N0_6_37 : std_logic;
	signal N0_6_38 : std_logic;
	signal N0_6_39 : std_logic;
	signal N0_6_40 : std_logic;
	signal N0_6_41 : std_logic;
	signal N0_6_42 : std_logic;
	signal N0_6_43 : std_logic;
	signal N0_6_44 : std_logic;
	signal N0_6_45 : std_logic;
	signal N0_6_46 : std_logic;
	signal N0_6_47 : std_logic;
	signal N0_6_48 : std_logic;
	signal N0_6_49 : std_logic;
	signal N0_6_50 : std_logic;
	signal N0_6_51 : std_logic;
	signal N0_6_52 : std_logic;
	signal N0_6_53 : std_logic;
	signal N0_6_54 : std_logic;
	signal N0_6_55 : std_logic;
	signal N0_6_56 : std_logic;
	signal N0_6_57 : std_logic;
	signal N0_6_58 : std_logic;
	signal N0_7_7 : std_logic;
	signal N0_7_8 : std_logic;
	signal N0_7_9 : std_logic;
	signal N0_7_10 : std_logic;
	signal N0_7_11 : std_logic;
	signal N0_7_12 : std_logic;
	signal N0_7_13 : std_logic;
	signal N0_7_14 : std_logic;
	signal N0_7_15 : std_logic;
	signal N0_7_16 : std_logic;
	signal N0_7_17 : std_logic;
	signal N0_7_18 : std_logic;
	signal N0_7_19 : std_logic;
	signal N0_7_20 : std_logic;
	signal N0_7_21 : std_logic;
	signal N0_7_22 : std_logic;
	signal N0_7_23 : std_logic;
	signal N0_7_24 : std_logic;
	signal N0_7_25 : std_logic;
	signal N0_7_26 : std_logic;
	signal N0_7_27 : std_logic;
	signal N0_7_28 : std_logic;
	signal N0_7_29 : std_logic;
	signal N0_7_30 : std_logic;
	signal N0_7_31 : std_logic;
	signal N0_7_32 : std_logic;
	signal N0_7_33 : std_logic;
	signal N0_7_34 : std_logic;
	signal N0_7_35 : std_logic;
	signal N0_7_36 : std_logic;
	signal N0_7_37 : std_logic;
	signal N0_7_38 : std_logic;
	signal N0_7_39 : std_logic;
	signal N0_7_40 : std_logic;
	signal N0_7_41 : std_logic;
	signal N0_7_42 : std_logic;
	signal N0_7_43 : std_logic;
	signal N0_7_44 : std_logic;
	signal N0_7_45 : std_logic;
	signal N0_7_46 : std_logic;
	signal N0_7_47 : std_logic;
	signal N0_7_48 : std_logic;
	signal N0_7_49 : std_logic;
	signal N0_7_50 : std_logic;
	signal N0_7_51 : std_logic;
	signal N0_7_52 : std_logic;
	signal N0_7_53 : std_logic;
	signal N0_7_54 : std_logic;
	signal N0_7_55 : std_logic;
	signal N0_7_56 : std_logic;
	signal N0_7_57 : std_logic;
	signal N0_7_58 : std_logic;
	signal N0_7_59 : std_logic;
	signal N0_8_8 : std_logic;
	signal N0_8_9 : std_logic;
	signal N0_8_10 : std_logic;
	signal N0_8_11 : std_logic;
	signal N0_8_12 : std_logic;
	signal N0_8_13 : std_logic;
	signal N0_8_14 : std_logic;
	signal N0_8_15 : std_logic;
	signal N0_8_16 : std_logic;
	signal N0_8_17 : std_logic;
	signal N0_8_18 : std_logic;
	signal N0_8_19 : std_logic;
	signal N0_8_20 : std_logic;
	signal N0_8_21 : std_logic;
	signal N0_8_22 : std_logic;
	signal N0_8_23 : std_logic;
	signal N0_8_24 : std_logic;
	signal N0_8_25 : std_logic;
	signal N0_8_26 : std_logic;
	signal N0_8_27 : std_logic;
	signal N0_8_28 : std_logic;
	signal N0_8_29 : std_logic;
	signal N0_8_30 : std_logic;
	signal N0_8_31 : std_logic;
	signal N0_8_32 : std_logic;
	signal N0_8_33 : std_logic;
	signal N0_8_34 : std_logic;
	signal N0_8_35 : std_logic;
	signal N0_8_36 : std_logic;
	signal N0_8_37 : std_logic;
	signal N0_8_38 : std_logic;
	signal N0_8_39 : std_logic;
	signal N0_8_40 : std_logic;
	signal N0_8_41 : std_logic;
	signal N0_8_42 : std_logic;
	signal N0_8_43 : std_logic;
	signal N0_8_44 : std_logic;
	signal N0_8_45 : std_logic;
	signal N0_8_46 : std_logic;
	signal N0_8_47 : std_logic;
	signal N0_8_48 : std_logic;
	signal N0_8_49 : std_logic;
	signal N0_8_50 : std_logic;
	signal N0_8_51 : std_logic;
	signal N0_8_52 : std_logic;
	signal N0_8_53 : std_logic;
	signal N0_8_54 : std_logic;
	signal N0_8_55 : std_logic;
	signal N0_8_56 : std_logic;
	signal N0_8_57 : std_logic;
	signal N0_8_58 : std_logic;
	signal N0_8_59 : std_logic;
	signal N0_8_60 : std_logic;
	signal N0_9_9 : std_logic;
	signal N0_9_10 : std_logic;
	signal N0_9_11 : std_logic;
	signal N0_9_12 : std_logic;
	signal N0_9_13 : std_logic;
	signal N0_9_14 : std_logic;
	signal N0_9_15 : std_logic;
	signal N0_9_16 : std_logic;
	signal N0_9_17 : std_logic;
	signal N0_9_18 : std_logic;
	signal N0_9_19 : std_logic;
	signal N0_9_20 : std_logic;
	signal N0_9_21 : std_logic;
	signal N0_9_22 : std_logic;
	signal N0_9_23 : std_logic;
	signal N0_9_24 : std_logic;
	signal N0_9_25 : std_logic;
	signal N0_9_26 : std_logic;
	signal N0_9_27 : std_logic;
	signal N0_9_28 : std_logic;
	signal N0_9_29 : std_logic;
	signal N0_9_30 : std_logic;
	signal N0_9_31 : std_logic;
	signal N0_9_32 : std_logic;
	signal N0_9_33 : std_logic;
	signal N0_9_34 : std_logic;
	signal N0_9_35 : std_logic;
	signal N0_9_36 : std_logic;
	signal N0_9_37 : std_logic;
	signal N0_9_38 : std_logic;
	signal N0_9_39 : std_logic;
	signal N0_9_40 : std_logic;
	signal N0_9_41 : std_logic;
	signal N0_9_42 : std_logic;
	signal N0_9_43 : std_logic;
	signal N0_9_44 : std_logic;
	signal N0_9_45 : std_logic;
	signal N0_9_46 : std_logic;
	signal N0_9_47 : std_logic;
	signal N0_9_48 : std_logic;
	signal N0_9_49 : std_logic;
	signal N0_9_50 : std_logic;
	signal N0_9_51 : std_logic;
	signal N0_9_52 : std_logic;
	signal N0_9_53 : std_logic;
	signal N0_9_54 : std_logic;
	signal N0_9_55 : std_logic;
	signal N0_9_56 : std_logic;
	signal N0_9_57 : std_logic;
	signal N0_9_58 : std_logic;
	signal N0_9_59 : std_logic;
	signal N0_9_60 : std_logic;
	signal N0_9_61 : std_logic;
	signal N0_10_10 : std_logic;
	signal N0_10_11 : std_logic;
	signal N0_10_12 : std_logic;
	signal N0_10_13 : std_logic;
	signal N0_10_14 : std_logic;
	signal N0_10_15 : std_logic;
	signal N0_10_16 : std_logic;
	signal N0_10_17 : std_logic;
	signal N0_10_18 : std_logic;
	signal N0_10_19 : std_logic;
	signal N0_10_20 : std_logic;
	signal N0_10_21 : std_logic;
	signal N0_10_22 : std_logic;
	signal N0_10_23 : std_logic;
	signal N0_10_24 : std_logic;
	signal N0_10_25 : std_logic;
	signal N0_10_26 : std_logic;
	signal N0_10_27 : std_logic;
	signal N0_10_28 : std_logic;
	signal N0_10_29 : std_logic;
	signal N0_10_30 : std_logic;
	signal N0_10_31 : std_logic;
	signal N0_10_32 : std_logic;
	signal N0_10_33 : std_logic;
	signal N0_10_34 : std_logic;
	signal N0_10_35 : std_logic;
	signal N0_10_36 : std_logic;
	signal N0_10_37 : std_logic;
	signal N0_10_38 : std_logic;
	signal N0_10_39 : std_logic;
	signal N0_10_40 : std_logic;
	signal N0_10_41 : std_logic;
	signal N0_10_42 : std_logic;
	signal N0_10_43 : std_logic;
	signal N0_10_44 : std_logic;
	signal N0_10_45 : std_logic;
	signal N0_10_46 : std_logic;
	signal N0_10_47 : std_logic;
	signal N0_10_48 : std_logic;
	signal N0_10_49 : std_logic;
	signal N0_10_50 : std_logic;
	signal N0_10_51 : std_logic;
	signal N0_10_52 : std_logic;
	signal N0_10_53 : std_logic;
	signal N0_10_54 : std_logic;
	signal N0_10_55 : std_logic;
	signal N0_10_56 : std_logic;
	signal N0_10_57 : std_logic;
	signal N0_10_58 : std_logic;
	signal N0_10_59 : std_logic;
	signal N0_10_60 : std_logic;
	signal N0_10_61 : std_logic;
	signal N0_10_62 : std_logic;
	signal N0_11_11 : std_logic;
	signal N0_11_12 : std_logic;
	signal N0_11_13 : std_logic;
	signal N0_11_14 : std_logic;
	signal N0_11_15 : std_logic;
	signal N0_11_16 : std_logic;
	signal N0_11_17 : std_logic;
	signal N0_11_18 : std_logic;
	signal N0_11_19 : std_logic;
	signal N0_11_20 : std_logic;
	signal N0_11_21 : std_logic;
	signal N0_11_22 : std_logic;
	signal N0_11_23 : std_logic;
	signal N0_11_24 : std_logic;
	signal N0_11_25 : std_logic;
	signal N0_11_26 : std_logic;
	signal N0_11_27 : std_logic;
	signal N0_11_28 : std_logic;
	signal N0_11_29 : std_logic;
	signal N0_11_30 : std_logic;
	signal N0_11_31 : std_logic;
	signal N0_11_32 : std_logic;
	signal N0_11_33 : std_logic;
	signal N0_11_34 : std_logic;
	signal N0_11_35 : std_logic;
	signal N0_11_36 : std_logic;
	signal N0_11_37 : std_logic;
	signal N0_11_38 : std_logic;
	signal N0_11_39 : std_logic;
	signal N0_11_40 : std_logic;
	signal N0_11_41 : std_logic;
	signal N0_11_42 : std_logic;
	signal N0_11_43 : std_logic;
	signal N0_11_44 : std_logic;
	signal N0_11_45 : std_logic;
	signal N0_11_46 : std_logic;
	signal N0_11_47 : std_logic;
	signal N0_11_48 : std_logic;
	signal N0_11_49 : std_logic;
	signal N0_11_50 : std_logic;
	signal N0_11_51 : std_logic;
	signal N0_11_52 : std_logic;
	signal N0_11_53 : std_logic;
	signal N0_11_54 : std_logic;
	signal N0_11_55 : std_logic;
	signal N0_11_56 : std_logic;
	signal N0_11_57 : std_logic;
	signal N0_11_58 : std_logic;
	signal N0_11_59 : std_logic;
	signal N0_11_60 : std_logic;
	signal N0_11_61 : std_logic;
	signal N0_11_62 : std_logic;
	signal N0_11_63 : std_logic;
	signal N0_12_12 : std_logic;
	signal N0_12_13 : std_logic;
	signal N0_12_14 : std_logic;
	signal N0_12_15 : std_logic;
	signal N0_12_16 : std_logic;
	signal N0_12_17 : std_logic;
	signal N0_12_18 : std_logic;
	signal N0_12_19 : std_logic;
	signal N0_12_20 : std_logic;
	signal N0_12_21 : std_logic;
	signal N0_12_22 : std_logic;
	signal N0_12_23 : std_logic;
	signal N0_12_24 : std_logic;
	signal N0_12_25 : std_logic;
	signal N0_12_26 : std_logic;
	signal N0_12_27 : std_logic;
	signal N0_12_28 : std_logic;
	signal N0_12_29 : std_logic;
	signal N0_12_30 : std_logic;
	signal N0_12_31 : std_logic;
	signal N0_12_32 : std_logic;
	signal N0_12_33 : std_logic;
	signal N0_12_34 : std_logic;
	signal N0_12_35 : std_logic;
	signal N0_12_36 : std_logic;
	signal N0_12_37 : std_logic;
	signal N0_12_38 : std_logic;
	signal N0_12_39 : std_logic;
	signal N0_12_40 : std_logic;
	signal N0_12_41 : std_logic;
	signal N0_12_42 : std_logic;
	signal N0_12_43 : std_logic;
	signal N0_12_44 : std_logic;
	signal N0_12_45 : std_logic;
	signal N0_12_46 : std_logic;
	signal N0_12_47 : std_logic;
	signal N0_12_48 : std_logic;
	signal N0_12_49 : std_logic;
	signal N0_12_50 : std_logic;
	signal N0_12_51 : std_logic;
	signal N0_12_52 : std_logic;
	signal N0_12_53 : std_logic;
	signal N0_12_54 : std_logic;
	signal N0_12_55 : std_logic;
	signal N0_12_56 : std_logic;
	signal N0_12_57 : std_logic;
	signal N0_12_58 : std_logic;
	signal N0_12_59 : std_logic;
	signal N0_12_60 : std_logic;
	signal N0_12_61 : std_logic;
	signal N0_12_62 : std_logic;
	signal N0_12_63 : std_logic;
	signal N0_12_64 : std_logic;
	signal N0_13_13 : std_logic;
	signal N0_13_14 : std_logic;
	signal N0_13_15 : std_logic;
	signal N0_13_16 : std_logic;
	signal N0_13_17 : std_logic;
	signal N0_13_18 : std_logic;
	signal N0_13_19 : std_logic;
	signal N0_13_20 : std_logic;
	signal N0_13_21 : std_logic;
	signal N0_13_22 : std_logic;
	signal N0_13_23 : std_logic;
	signal N0_13_24 : std_logic;
	signal N0_13_25 : std_logic;
	signal N0_13_26 : std_logic;
	signal N0_13_27 : std_logic;
	signal N0_13_28 : std_logic;
	signal N0_13_29 : std_logic;
	signal N0_13_30 : std_logic;
	signal N0_13_31 : std_logic;
	signal N0_13_32 : std_logic;
	signal N0_13_33 : std_logic;
	signal N0_13_34 : std_logic;
	signal N0_13_35 : std_logic;
	signal N0_13_36 : std_logic;
	signal N0_13_37 : std_logic;
	signal N0_13_38 : std_logic;
	signal N0_13_39 : std_logic;
	signal N0_13_40 : std_logic;
	signal N0_13_41 : std_logic;
	signal N0_13_42 : std_logic;
	signal N0_13_43 : std_logic;
	signal N0_13_44 : std_logic;
	signal N0_13_45 : std_logic;
	signal N0_13_46 : std_logic;
	signal N0_13_47 : std_logic;
	signal N0_13_48 : std_logic;
	signal N0_13_49 : std_logic;
	signal N0_13_50 : std_logic;
	signal N0_13_51 : std_logic;
	signal N0_13_52 : std_logic;
	signal N0_13_53 : std_logic;
	signal N0_13_54 : std_logic;
	signal N0_13_55 : std_logic;
	signal N0_13_56 : std_logic;
	signal N0_13_57 : std_logic;
	signal N0_13_58 : std_logic;
	signal N0_13_59 : std_logic;
	signal N0_13_60 : std_logic;
	signal N0_13_61 : std_logic;
	signal N0_13_62 : std_logic;
	signal N0_13_63 : std_logic;
	signal N0_13_64 : std_logic;
	signal N0_13_65 : std_logic;
	signal N0_14_14 : std_logic;
	signal N0_14_15 : std_logic;
	signal N0_14_16 : std_logic;
	signal N0_14_17 : std_logic;
	signal N0_14_18 : std_logic;
	signal N0_14_19 : std_logic;
	signal N0_14_20 : std_logic;
	signal N0_14_21 : std_logic;
	signal N0_14_22 : std_logic;
	signal N0_14_23 : std_logic;
	signal N0_14_24 : std_logic;
	signal N0_14_25 : std_logic;
	signal N0_14_26 : std_logic;
	signal N0_14_27 : std_logic;
	signal N0_14_28 : std_logic;
	signal N0_14_29 : std_logic;
	signal N0_14_30 : std_logic;
	signal N0_14_31 : std_logic;
	signal N0_14_32 : std_logic;
	signal N0_14_33 : std_logic;
	signal N0_14_34 : std_logic;
	signal N0_14_35 : std_logic;
	signal N0_14_36 : std_logic;
	signal N0_14_37 : std_logic;
	signal N0_14_38 : std_logic;
	signal N0_14_39 : std_logic;
	signal N0_14_40 : std_logic;
	signal N0_14_41 : std_logic;
	signal N0_14_42 : std_logic;
	signal N0_14_43 : std_logic;
	signal N0_14_44 : std_logic;
	signal N0_14_45 : std_logic;
	signal N0_14_46 : std_logic;
	signal N0_14_47 : std_logic;
	signal N0_14_48 : std_logic;
	signal N0_14_49 : std_logic;
	signal N0_14_50 : std_logic;
	signal N0_14_51 : std_logic;
	signal N0_14_52 : std_logic;
	signal N0_14_53 : std_logic;
	signal N0_14_54 : std_logic;
	signal N0_14_55 : std_logic;
	signal N0_14_56 : std_logic;
	signal N0_14_57 : std_logic;
	signal N0_14_58 : std_logic;
	signal N0_14_59 : std_logic;
	signal N0_14_60 : std_logic;
	signal N0_14_61 : std_logic;
	signal N0_14_62 : std_logic;
	signal N0_14_63 : std_logic;
	signal N0_14_64 : std_logic;
	signal N0_14_65 : std_logic;
	signal N0_14_66 : std_logic;
	signal N0_15_15 : std_logic;
	signal N0_15_16 : std_logic;
	signal N0_15_17 : std_logic;
	signal N0_15_18 : std_logic;
	signal N0_15_19 : std_logic;
	signal N0_15_20 : std_logic;
	signal N0_15_21 : std_logic;
	signal N0_15_22 : std_logic;
	signal N0_15_23 : std_logic;
	signal N0_15_24 : std_logic;
	signal N0_15_25 : std_logic;
	signal N0_15_26 : std_logic;
	signal N0_15_27 : std_logic;
	signal N0_15_28 : std_logic;
	signal N0_15_29 : std_logic;
	signal N0_15_30 : std_logic;
	signal N0_15_31 : std_logic;
	signal N0_15_32 : std_logic;
	signal N0_15_33 : std_logic;
	signal N0_15_34 : std_logic;
	signal N0_15_35 : std_logic;
	signal N0_15_36 : std_logic;
	signal N0_15_37 : std_logic;
	signal N0_15_38 : std_logic;
	signal N0_15_39 : std_logic;
	signal N0_15_40 : std_logic;
	signal N0_15_41 : std_logic;
	signal N0_15_42 : std_logic;
	signal N0_15_43 : std_logic;
	signal N0_15_44 : std_logic;
	signal N0_15_45 : std_logic;
	signal N0_15_46 : std_logic;
	signal N0_15_47 : std_logic;
	signal N0_15_48 : std_logic;
	signal N0_15_49 : std_logic;
	signal N0_15_50 : std_logic;
	signal N0_15_51 : std_logic;
	signal N0_15_52 : std_logic;
	signal N0_15_53 : std_logic;
	signal N0_15_54 : std_logic;
	signal N0_15_55 : std_logic;
	signal N0_15_56 : std_logic;
	signal N0_15_57 : std_logic;
	signal N0_15_58 : std_logic;
	signal N0_15_59 : std_logic;
	signal N0_15_60 : std_logic;
	signal N0_15_61 : std_logic;
	signal N0_15_62 : std_logic;
	signal N0_15_63 : std_logic;
	signal N0_15_64 : std_logic;
	signal N0_15_65 : std_logic;
	signal N0_15_66 : std_logic;
	signal N0_15_67 : std_logic;
	signal N0_16_16 : std_logic;
	signal N0_16_17 : std_logic;
	signal N0_16_18 : std_logic;
	signal N0_16_19 : std_logic;
	signal N0_16_20 : std_logic;
	signal N0_16_21 : std_logic;
	signal N0_16_22 : std_logic;
	signal N0_16_23 : std_logic;
	signal N0_16_24 : std_logic;
	signal N0_16_25 : std_logic;
	signal N0_16_26 : std_logic;
	signal N0_16_27 : std_logic;
	signal N0_16_28 : std_logic;
	signal N0_16_29 : std_logic;
	signal N0_16_30 : std_logic;
	signal N0_16_31 : std_logic;
	signal N0_16_32 : std_logic;
	signal N0_16_33 : std_logic;
	signal N0_16_34 : std_logic;
	signal N0_16_35 : std_logic;
	signal N0_16_36 : std_logic;
	signal N0_16_37 : std_logic;
	signal N0_16_38 : std_logic;
	signal N0_16_39 : std_logic;
	signal N0_16_40 : std_logic;
	signal N0_16_41 : std_logic;
	signal N0_16_42 : std_logic;
	signal N0_16_43 : std_logic;
	signal N0_16_44 : std_logic;
	signal N0_16_45 : std_logic;
	signal N0_16_46 : std_logic;
	signal N0_16_47 : std_logic;
	signal N0_16_48 : std_logic;
	signal N0_16_49 : std_logic;
	signal N0_16_50 : std_logic;
	signal N0_16_51 : std_logic;
	signal N0_16_52 : std_logic;
	signal N0_16_53 : std_logic;
	signal N0_16_54 : std_logic;
	signal N0_16_55 : std_logic;
	signal N0_16_56 : std_logic;
	signal N0_16_57 : std_logic;
	signal N0_16_58 : std_logic;
	signal N0_16_59 : std_logic;
	signal N0_16_60 : std_logic;
	signal N0_16_61 : std_logic;
	signal N0_16_62 : std_logic;
	signal N0_16_63 : std_logic;
	signal N0_16_64 : std_logic;
	signal N0_16_65 : std_logic;
	signal N0_16_66 : std_logic;
	signal N0_16_67 : std_logic;
	signal N0_16_68 : std_logic;
	signal N0_17_17 : std_logic;
	signal N0_17_18 : std_logic;
	signal N0_17_19 : std_logic;
	signal N0_17_20 : std_logic;
	signal N0_17_21 : std_logic;
	signal N0_17_22 : std_logic;
	signal N0_17_23 : std_logic;
	signal N0_17_24 : std_logic;
	signal N0_17_25 : std_logic;
	signal N0_17_26 : std_logic;
	signal N0_17_27 : std_logic;
	signal N0_17_28 : std_logic;
	signal N0_17_29 : std_logic;
	signal N0_17_30 : std_logic;
	signal N0_17_31 : std_logic;
	signal N0_17_32 : std_logic;
	signal N0_17_33 : std_logic;
	signal N0_17_34 : std_logic;
	signal N0_17_35 : std_logic;
	signal N0_17_36 : std_logic;
	signal N0_17_37 : std_logic;
	signal N0_17_38 : std_logic;
	signal N0_17_39 : std_logic;
	signal N0_17_40 : std_logic;
	signal N0_17_41 : std_logic;
	signal N0_17_42 : std_logic;
	signal N0_17_43 : std_logic;
	signal N0_17_44 : std_logic;
	signal N0_17_45 : std_logic;
	signal N0_17_46 : std_logic;
	signal N0_17_47 : std_logic;
	signal N0_17_48 : std_logic;
	signal N0_17_49 : std_logic;
	signal N0_17_50 : std_logic;
	signal N0_17_51 : std_logic;
	signal N0_17_52 : std_logic;
	signal N0_17_53 : std_logic;
	signal N0_17_54 : std_logic;
	signal N0_17_55 : std_logic;
	signal N0_17_56 : std_logic;
	signal N0_17_57 : std_logic;
	signal N0_17_58 : std_logic;
	signal N0_17_59 : std_logic;
	signal N0_17_60 : std_logic;
	signal N0_17_61 : std_logic;
	signal N0_17_62 : std_logic;
	signal N0_17_63 : std_logic;
	signal N0_17_64 : std_logic;
	signal N0_17_65 : std_logic;
	signal N0_17_66 : std_logic;
	signal N0_17_67 : std_logic;
	signal N0_17_68 : std_logic;
	signal N0_17_69 : std_logic;
	signal N0_18_18 : std_logic;
	signal N0_18_19 : std_logic;
	signal N0_18_20 : std_logic;
	signal N0_18_21 : std_logic;
	signal N0_18_22 : std_logic;
	signal N0_18_23 : std_logic;
	signal N0_18_24 : std_logic;
	signal N0_18_25 : std_logic;
	signal N0_18_26 : std_logic;
	signal N0_18_27 : std_logic;
	signal N0_18_28 : std_logic;
	signal N0_18_29 : std_logic;
	signal N0_18_30 : std_logic;
	signal N0_18_31 : std_logic;
	signal N0_18_32 : std_logic;
	signal N0_18_33 : std_logic;
	signal N0_18_34 : std_logic;
	signal N0_18_35 : std_logic;
	signal N0_18_36 : std_logic;
	signal N0_18_37 : std_logic;
	signal N0_18_38 : std_logic;
	signal N0_18_39 : std_logic;
	signal N0_18_40 : std_logic;
	signal N0_18_41 : std_logic;
	signal N0_18_42 : std_logic;
	signal N0_18_43 : std_logic;
	signal N0_18_44 : std_logic;
	signal N0_18_45 : std_logic;
	signal N0_18_46 : std_logic;
	signal N0_18_47 : std_logic;
	signal N0_18_48 : std_logic;
	signal N0_18_49 : std_logic;
	signal N0_18_50 : std_logic;
	signal N0_18_51 : std_logic;
	signal N0_18_52 : std_logic;
	signal N0_18_53 : std_logic;
	signal N0_18_54 : std_logic;
	signal N0_18_55 : std_logic;
	signal N0_18_56 : std_logic;
	signal N0_18_57 : std_logic;
	signal N0_18_58 : std_logic;
	signal N0_18_59 : std_logic;
	signal N0_18_60 : std_logic;
	signal N0_18_61 : std_logic;
	signal N0_18_62 : std_logic;
	signal N0_18_63 : std_logic;
	signal N0_18_64 : std_logic;
	signal N0_18_65 : std_logic;
	signal N0_18_66 : std_logic;
	signal N0_18_67 : std_logic;
	signal N0_18_68 : std_logic;
	signal N0_18_69 : std_logic;
	signal N0_18_70 : std_logic;
	signal N0_19_19 : std_logic;
	signal N0_19_20 : std_logic;
	signal N0_19_21 : std_logic;
	signal N0_19_22 : std_logic;
	signal N0_19_23 : std_logic;
	signal N0_19_24 : std_logic;
	signal N0_19_25 : std_logic;
	signal N0_19_26 : std_logic;
	signal N0_19_27 : std_logic;
	signal N0_19_28 : std_logic;
	signal N0_19_29 : std_logic;
	signal N0_19_30 : std_logic;
	signal N0_19_31 : std_logic;
	signal N0_19_32 : std_logic;
	signal N0_19_33 : std_logic;
	signal N0_19_34 : std_logic;
	signal N0_19_35 : std_logic;
	signal N0_19_36 : std_logic;
	signal N0_19_37 : std_logic;
	signal N0_19_38 : std_logic;
	signal N0_19_39 : std_logic;
	signal N0_19_40 : std_logic;
	signal N0_19_41 : std_logic;
	signal N0_19_42 : std_logic;
	signal N0_19_43 : std_logic;
	signal N0_19_44 : std_logic;
	signal N0_19_45 : std_logic;
	signal N0_19_46 : std_logic;
	signal N0_19_47 : std_logic;
	signal N0_19_48 : std_logic;
	signal N0_19_49 : std_logic;
	signal N0_19_50 : std_logic;
	signal N0_19_51 : std_logic;
	signal N0_19_52 : std_logic;
	signal N0_19_53 : std_logic;
	signal N0_19_54 : std_logic;
	signal N0_19_55 : std_logic;
	signal N0_19_56 : std_logic;
	signal N0_19_57 : std_logic;
	signal N0_19_58 : std_logic;
	signal N0_19_59 : std_logic;
	signal N0_19_60 : std_logic;
	signal N0_19_61 : std_logic;
	signal N0_19_62 : std_logic;
	signal N0_19_63 : std_logic;
	signal N0_19_64 : std_logic;
	signal N0_19_65 : std_logic;
	signal N0_19_66 : std_logic;
	signal N0_19_67 : std_logic;
	signal N0_19_68 : std_logic;
	signal N0_19_69 : std_logic;
	signal N0_19_70 : std_logic;
	signal N0_19_71 : std_logic;
	signal N0_20_20 : std_logic;
	signal N0_20_21 : std_logic;
	signal N0_20_22 : std_logic;
	signal N0_20_23 : std_logic;
	signal N0_20_24 : std_logic;
	signal N0_20_25 : std_logic;
	signal N0_20_26 : std_logic;
	signal N0_20_27 : std_logic;
	signal N0_20_28 : std_logic;
	signal N0_20_29 : std_logic;
	signal N0_20_30 : std_logic;
	signal N0_20_31 : std_logic;
	signal N0_20_32 : std_logic;
	signal N0_20_33 : std_logic;
	signal N0_20_34 : std_logic;
	signal N0_20_35 : std_logic;
	signal N0_20_36 : std_logic;
	signal N0_20_37 : std_logic;
	signal N0_20_38 : std_logic;
	signal N0_20_39 : std_logic;
	signal N0_20_40 : std_logic;
	signal N0_20_41 : std_logic;
	signal N0_20_42 : std_logic;
	signal N0_20_43 : std_logic;
	signal N0_20_44 : std_logic;
	signal N0_20_45 : std_logic;
	signal N0_20_46 : std_logic;
	signal N0_20_47 : std_logic;
	signal N0_20_48 : std_logic;
	signal N0_20_49 : std_logic;
	signal N0_20_50 : std_logic;
	signal N0_20_51 : std_logic;
	signal N0_20_52 : std_logic;
	signal N0_20_53 : std_logic;
	signal N0_20_54 : std_logic;
	signal N0_20_55 : std_logic;
	signal N0_20_56 : std_logic;
	signal N0_20_57 : std_logic;
	signal N0_20_58 : std_logic;
	signal N0_20_59 : std_logic;
	signal N0_20_60 : std_logic;
	signal N0_20_61 : std_logic;
	signal N0_20_62 : std_logic;
	signal N0_20_63 : std_logic;
	signal N0_20_64 : std_logic;
	signal N0_20_65 : std_logic;
	signal N0_20_66 : std_logic;
	signal N0_20_67 : std_logic;
	signal N0_20_68 : std_logic;
	signal N0_20_69 : std_logic;
	signal N0_20_70 : std_logic;
	signal N0_20_71 : std_logic;
	signal N0_20_72 : std_logic;
	signal N0_21_21 : std_logic;
	signal N0_21_22 : std_logic;
	signal N0_21_23 : std_logic;
	signal N0_21_24 : std_logic;
	signal N0_21_25 : std_logic;
	signal N0_21_26 : std_logic;
	signal N0_21_27 : std_logic;
	signal N0_21_28 : std_logic;
	signal N0_21_29 : std_logic;
	signal N0_21_30 : std_logic;
	signal N0_21_31 : std_logic;
	signal N0_21_32 : std_logic;
	signal N0_21_33 : std_logic;
	signal N0_21_34 : std_logic;
	signal N0_21_35 : std_logic;
	signal N0_21_36 : std_logic;
	signal N0_21_37 : std_logic;
	signal N0_21_38 : std_logic;
	signal N0_21_39 : std_logic;
	signal N0_21_40 : std_logic;
	signal N0_21_41 : std_logic;
	signal N0_21_42 : std_logic;
	signal N0_21_43 : std_logic;
	signal N0_21_44 : std_logic;
	signal N0_21_45 : std_logic;
	signal N0_21_46 : std_logic;
	signal N0_21_47 : std_logic;
	signal N0_21_48 : std_logic;
	signal N0_21_49 : std_logic;
	signal N0_21_50 : std_logic;
	signal N0_21_51 : std_logic;
	signal N0_21_52 : std_logic;
	signal N0_21_53 : std_logic;
	signal N0_21_54 : std_logic;
	signal N0_21_55 : std_logic;
	signal N0_21_56 : std_logic;
	signal N0_21_57 : std_logic;
	signal N0_21_58 : std_logic;
	signal N0_21_59 : std_logic;
	signal N0_21_60 : std_logic;
	signal N0_21_61 : std_logic;
	signal N0_21_62 : std_logic;
	signal N0_21_63 : std_logic;
	signal N0_21_64 : std_logic;
	signal N0_21_65 : std_logic;
	signal N0_21_66 : std_logic;
	signal N0_21_67 : std_logic;
	signal N0_21_68 : std_logic;
	signal N0_21_69 : std_logic;
	signal N0_21_70 : std_logic;
	signal N0_21_71 : std_logic;
	signal N0_21_72 : std_logic;
	signal N0_21_73 : std_logic;
	signal N0_22_22 : std_logic;
	signal N0_22_23 : std_logic;
	signal N0_22_24 : std_logic;
	signal N0_22_25 : std_logic;
	signal N0_22_26 : std_logic;
	signal N0_22_27 : std_logic;
	signal N0_22_28 : std_logic;
	signal N0_22_29 : std_logic;
	signal N0_22_30 : std_logic;
	signal N0_22_31 : std_logic;
	signal N0_22_32 : std_logic;
	signal N0_22_33 : std_logic;
	signal N0_22_34 : std_logic;
	signal N0_22_35 : std_logic;
	signal N0_22_36 : std_logic;
	signal N0_22_37 : std_logic;
	signal N0_22_38 : std_logic;
	signal N0_22_39 : std_logic;
	signal N0_22_40 : std_logic;
	signal N0_22_41 : std_logic;
	signal N0_22_42 : std_logic;
	signal N0_22_43 : std_logic;
	signal N0_22_44 : std_logic;
	signal N0_22_45 : std_logic;
	signal N0_22_46 : std_logic;
	signal N0_22_47 : std_logic;
	signal N0_22_48 : std_logic;
	signal N0_22_49 : std_logic;
	signal N0_22_50 : std_logic;
	signal N0_22_51 : std_logic;
	signal N0_22_52 : std_logic;
	signal N0_22_53 : std_logic;
	signal N0_22_54 : std_logic;
	signal N0_22_55 : std_logic;
	signal N0_22_56 : std_logic;
	signal N0_22_57 : std_logic;
	signal N0_22_58 : std_logic;
	signal N0_22_59 : std_logic;
	signal N0_22_60 : std_logic;
	signal N0_22_61 : std_logic;
	signal N0_22_62 : std_logic;
	signal N0_22_63 : std_logic;
	signal N0_22_64 : std_logic;
	signal N0_22_65 : std_logic;
	signal N0_22_66 : std_logic;
	signal N0_22_67 : std_logic;
	signal N0_22_68 : std_logic;
	signal N0_22_69 : std_logic;
	signal N0_22_70 : std_logic;
	signal N0_22_71 : std_logic;
	signal N0_22_72 : std_logic;
	signal N0_22_73 : std_logic;
	signal N0_22_74 : std_logic;
	signal N0_23_23 : std_logic;
	signal N0_23_24 : std_logic;
	signal N0_23_25 : std_logic;
	signal N0_23_26 : std_logic;
	signal N0_23_27 : std_logic;
	signal N0_23_28 : std_logic;
	signal N0_23_29 : std_logic;
	signal N0_23_30 : std_logic;
	signal N0_23_31 : std_logic;
	signal N0_23_32 : std_logic;
	signal N0_23_33 : std_logic;
	signal N0_23_34 : std_logic;
	signal N0_23_35 : std_logic;
	signal N0_23_36 : std_logic;
	signal N0_23_37 : std_logic;
	signal N0_23_38 : std_logic;
	signal N0_23_39 : std_logic;
	signal N0_23_40 : std_logic;
	signal N0_23_41 : std_logic;
	signal N0_23_42 : std_logic;
	signal N0_23_43 : std_logic;
	signal N0_23_44 : std_logic;
	signal N0_23_45 : std_logic;
	signal N0_23_46 : std_logic;
	signal N0_23_47 : std_logic;
	signal N0_23_48 : std_logic;
	signal N0_23_49 : std_logic;
	signal N0_23_50 : std_logic;
	signal N0_23_51 : std_logic;
	signal N0_23_52 : std_logic;
	signal N0_23_53 : std_logic;
	signal N0_23_54 : std_logic;
	signal N0_23_55 : std_logic;
	signal N0_23_56 : std_logic;
	signal N0_23_57 : std_logic;
	signal N0_23_58 : std_logic;
	signal N0_23_59 : std_logic;
	signal N0_23_60 : std_logic;
	signal N0_23_61 : std_logic;
	signal N0_23_62 : std_logic;
	signal N0_23_63 : std_logic;
	signal N0_23_64 : std_logic;
	signal N0_23_65 : std_logic;
	signal N0_23_66 : std_logic;
	signal N0_23_67 : std_logic;
	signal N0_23_68 : std_logic;
	signal N0_23_69 : std_logic;
	signal N0_23_70 : std_logic;
	signal N0_23_71 : std_logic;
	signal N0_23_72 : std_logic;
	signal N0_23_73 : std_logic;
	signal N0_23_74 : std_logic;
	signal N0_23_75 : std_logic;
	signal N0_24_24 : std_logic;
	signal N0_24_25 : std_logic;
	signal N0_24_26 : std_logic;
	signal N0_24_27 : std_logic;
	signal N0_24_28 : std_logic;
	signal N0_24_29 : std_logic;
	signal N0_24_30 : std_logic;
	signal N0_24_31 : std_logic;
	signal N0_24_32 : std_logic;
	signal N0_24_33 : std_logic;
	signal N0_24_34 : std_logic;
	signal N0_24_35 : std_logic;
	signal N0_24_36 : std_logic;
	signal N0_24_37 : std_logic;
	signal N0_24_38 : std_logic;
	signal N0_24_39 : std_logic;
	signal N0_24_40 : std_logic;
	signal N0_24_41 : std_logic;
	signal N0_24_42 : std_logic;
	signal N0_24_43 : std_logic;
	signal N0_24_44 : std_logic;
	signal N0_24_45 : std_logic;
	signal N0_24_46 : std_logic;
	signal N0_24_47 : std_logic;
	signal N0_24_48 : std_logic;
	signal N0_24_49 : std_logic;
	signal N0_24_50 : std_logic;
	signal N0_24_51 : std_logic;
	signal N0_24_52 : std_logic;
	signal N0_24_53 : std_logic;
	signal N0_24_54 : std_logic;
	signal N0_24_55 : std_logic;
	signal N0_24_56 : std_logic;
	signal N0_24_57 : std_logic;
	signal N0_24_58 : std_logic;
	signal N0_24_59 : std_logic;
	signal N0_24_60 : std_logic;
	signal N0_24_61 : std_logic;
	signal N0_24_62 : std_logic;
	signal N0_24_63 : std_logic;
	signal N0_24_64 : std_logic;
	signal N0_24_65 : std_logic;
	signal N0_24_66 : std_logic;
	signal N0_24_67 : std_logic;
	signal N0_24_68 : std_logic;
	signal N0_24_69 : std_logic;
	signal N0_24_70 : std_logic;
	signal N0_24_71 : std_logic;
	signal N0_24_72 : std_logic;
	signal N0_24_73 : std_logic;
	signal N0_24_74 : std_logic;
	signal N0_24_75 : std_logic;
	signal N0_24_76 : std_logic;
	signal N0_25_25 : std_logic;
	signal N0_25_26 : std_logic;
	signal N0_25_27 : std_logic;
	signal N0_25_28 : std_logic;
	signal N0_25_29 : std_logic;
	signal N0_25_30 : std_logic;
	signal N0_25_31 : std_logic;
	signal N0_25_32 : std_logic;
	signal N0_25_33 : std_logic;
	signal N0_25_34 : std_logic;
	signal N0_25_35 : std_logic;
	signal N0_25_36 : std_logic;
	signal N0_25_37 : std_logic;
	signal N0_25_38 : std_logic;
	signal N0_25_39 : std_logic;
	signal N0_25_40 : std_logic;
	signal N0_25_41 : std_logic;
	signal N0_25_42 : std_logic;
	signal N0_25_43 : std_logic;
	signal N0_25_44 : std_logic;
	signal N0_25_45 : std_logic;
	signal N0_25_46 : std_logic;
	signal N0_25_47 : std_logic;
	signal N0_25_48 : std_logic;
	signal N0_25_49 : std_logic;
	signal N0_25_50 : std_logic;
	signal N0_25_51 : std_logic;
	signal N0_25_52 : std_logic;
	signal N0_25_53 : std_logic;
	signal N0_25_54 : std_logic;
	signal N0_25_55 : std_logic;
	signal N0_25_56 : std_logic;
	signal N0_25_57 : std_logic;
	signal N0_25_58 : std_logic;
	signal N0_25_59 : std_logic;
	signal N0_25_60 : std_logic;
	signal N0_25_61 : std_logic;
	signal N0_25_62 : std_logic;
	signal N0_25_63 : std_logic;
	signal N0_25_64 : std_logic;
	signal N0_25_65 : std_logic;
	signal N0_25_66 : std_logic;
	signal N0_25_67 : std_logic;
	signal N0_25_68 : std_logic;
	signal N0_25_69 : std_logic;
	signal N0_25_70 : std_logic;
	signal N0_25_71 : std_logic;
	signal N0_25_72 : std_logic;
	signal N0_25_73 : std_logic;
	signal N0_25_74 : std_logic;
	signal N0_25_75 : std_logic;
	signal N0_25_76 : std_logic;
	signal N0_25_77 : std_logic;
	signal N0_26_26 : std_logic;
	signal N0_26_27 : std_logic;
	signal N0_26_28 : std_logic;
	signal N0_26_29 : std_logic;
	signal N0_26_30 : std_logic;
	signal N0_26_31 : std_logic;
	signal N0_26_32 : std_logic;
	signal N0_26_33 : std_logic;
	signal N0_26_34 : std_logic;
	signal N0_26_35 : std_logic;
	signal N0_26_36 : std_logic;
	signal N0_26_37 : std_logic;
	signal N0_26_38 : std_logic;
	signal N0_26_39 : std_logic;
	signal N0_26_40 : std_logic;
	signal N0_26_41 : std_logic;
	signal N0_26_42 : std_logic;
	signal N0_26_43 : std_logic;
	signal N0_26_44 : std_logic;
	signal N0_26_45 : std_logic;
	signal N0_26_46 : std_logic;
	signal N0_26_47 : std_logic;
	signal N0_26_48 : std_logic;
	signal N0_26_49 : std_logic;
	signal N0_26_50 : std_logic;
	signal N0_26_51 : std_logic;
	signal N0_26_52 : std_logic;
	signal N0_26_53 : std_logic;
	signal N0_26_54 : std_logic;
	signal N0_26_55 : std_logic;
	signal N0_26_56 : std_logic;
	signal N0_26_57 : std_logic;
	signal N0_26_58 : std_logic;
	signal N0_26_59 : std_logic;
	signal N0_26_60 : std_logic;
	signal N0_26_61 : std_logic;
	signal N0_26_62 : std_logic;
	signal N0_26_63 : std_logic;
	signal N0_26_64 : std_logic;
	signal N0_26_65 : std_logic;
	signal N0_26_66 : std_logic;
	signal N0_26_67 : std_logic;
	signal N0_26_68 : std_logic;
	signal N0_26_69 : std_logic;
	signal N0_26_70 : std_logic;
	signal N0_26_71 : std_logic;
	signal N0_26_72 : std_logic;
	signal N0_26_73 : std_logic;
	signal N0_26_74 : std_logic;
	signal N0_26_75 : std_logic;
	signal N0_26_76 : std_logic;
	signal N0_26_77 : std_logic;
	signal N0_26_78 : std_logic;
	signal N0_27_27 : std_logic;
	signal N0_27_28 : std_logic;
	signal N0_27_29 : std_logic;
	signal N0_27_30 : std_logic;
	signal N0_27_31 : std_logic;
	signal N0_27_32 : std_logic;
	signal N0_27_33 : std_logic;
	signal N0_27_34 : std_logic;
	signal N0_27_35 : std_logic;
	signal N0_27_36 : std_logic;
	signal N0_27_37 : std_logic;
	signal N0_27_38 : std_logic;
	signal N0_27_39 : std_logic;
	signal N0_27_40 : std_logic;
	signal N0_27_41 : std_logic;
	signal N0_27_42 : std_logic;
	signal N0_27_43 : std_logic;
	signal N0_27_44 : std_logic;
	signal N0_27_45 : std_logic;
	signal N0_27_46 : std_logic;
	signal N0_27_47 : std_logic;
	signal N0_27_48 : std_logic;
	signal N0_27_49 : std_logic;
	signal N0_27_50 : std_logic;
	signal N0_27_51 : std_logic;
	signal N0_27_52 : std_logic;
	signal N0_27_53 : std_logic;
	signal N0_27_54 : std_logic;
	signal N0_27_55 : std_logic;
	signal N0_27_56 : std_logic;
	signal N0_27_57 : std_logic;
	signal N0_27_58 : std_logic;
	signal N0_27_59 : std_logic;
	signal N0_27_60 : std_logic;
	signal N0_27_61 : std_logic;
	signal N0_27_62 : std_logic;
	signal N0_27_63 : std_logic;
	signal N0_27_64 : std_logic;
	signal N0_27_65 : std_logic;
	signal N0_27_66 : std_logic;
	signal N0_27_67 : std_logic;
	signal N0_27_68 : std_logic;
	signal N0_27_69 : std_logic;
	signal N0_27_70 : std_logic;
	signal N0_27_71 : std_logic;
	signal N0_27_72 : std_logic;
	signal N0_27_73 : std_logic;
	signal N0_27_74 : std_logic;
	signal N0_27_75 : std_logic;
	signal N0_27_76 : std_logic;
	signal N0_27_77 : std_logic;
	signal N0_27_78 : std_logic;
	signal N0_27_79 : std_logic;
	signal N0_28_28 : std_logic;
	signal N0_28_29 : std_logic;
	signal N0_28_30 : std_logic;
	signal N0_28_31 : std_logic;
	signal N0_28_32 : std_logic;
	signal N0_28_33 : std_logic;
	signal N0_28_34 : std_logic;
	signal N0_28_35 : std_logic;
	signal N0_28_36 : std_logic;
	signal N0_28_37 : std_logic;
	signal N0_28_38 : std_logic;
	signal N0_28_39 : std_logic;
	signal N0_28_40 : std_logic;
	signal N0_28_41 : std_logic;
	signal N0_28_42 : std_logic;
	signal N0_28_43 : std_logic;
	signal N0_28_44 : std_logic;
	signal N0_28_45 : std_logic;
	signal N0_28_46 : std_logic;
	signal N0_28_47 : std_logic;
	signal N0_28_48 : std_logic;
	signal N0_28_49 : std_logic;
	signal N0_28_50 : std_logic;
	signal N0_28_51 : std_logic;
	signal N0_28_52 : std_logic;
	signal N0_28_53 : std_logic;
	signal N0_28_54 : std_logic;
	signal N0_28_55 : std_logic;
	signal N0_28_56 : std_logic;
	signal N0_28_57 : std_logic;
	signal N0_28_58 : std_logic;
	signal N0_28_59 : std_logic;
	signal N0_28_60 : std_logic;
	signal N0_28_61 : std_logic;
	signal N0_28_62 : std_logic;
	signal N0_28_63 : std_logic;
	signal N0_28_64 : std_logic;
	signal N0_28_65 : std_logic;
	signal N0_28_66 : std_logic;
	signal N0_28_67 : std_logic;
	signal N0_28_68 : std_logic;
	signal N0_28_69 : std_logic;
	signal N0_28_70 : std_logic;
	signal N0_28_71 : std_logic;
	signal N0_28_72 : std_logic;
	signal N0_28_73 : std_logic;
	signal N0_28_74 : std_logic;
	signal N0_28_75 : std_logic;
	signal N0_28_76 : std_logic;
	signal N0_28_77 : std_logic;
	signal N0_28_78 : std_logic;
	signal N0_28_79 : std_logic;
	signal N0_28_80 : std_logic;
	signal N0_29_29 : std_logic;
	signal N0_29_30 : std_logic;
	signal N0_29_31 : std_logic;
	signal N0_29_32 : std_logic;
	signal N0_29_33 : std_logic;
	signal N0_29_34 : std_logic;
	signal N0_29_35 : std_logic;
	signal N0_29_36 : std_logic;
	signal N0_29_37 : std_logic;
	signal N0_29_38 : std_logic;
	signal N0_29_39 : std_logic;
	signal N0_29_40 : std_logic;
	signal N0_29_41 : std_logic;
	signal N0_29_42 : std_logic;
	signal N0_29_43 : std_logic;
	signal N0_29_44 : std_logic;
	signal N0_29_45 : std_logic;
	signal N0_29_46 : std_logic;
	signal N0_29_47 : std_logic;
	signal N0_29_48 : std_logic;
	signal N0_29_49 : std_logic;
	signal N0_29_50 : std_logic;
	signal N0_29_51 : std_logic;
	signal N0_29_52 : std_logic;
	signal N0_29_53 : std_logic;
	signal N0_29_54 : std_logic;
	signal N0_29_55 : std_logic;
	signal N0_29_56 : std_logic;
	signal N0_29_57 : std_logic;
	signal N0_29_58 : std_logic;
	signal N0_29_59 : std_logic;
	signal N0_29_60 : std_logic;
	signal N0_29_61 : std_logic;
	signal N0_29_62 : std_logic;
	signal N0_29_63 : std_logic;
	signal N0_29_64 : std_logic;
	signal N0_29_65 : std_logic;
	signal N0_29_66 : std_logic;
	signal N0_29_67 : std_logic;
	signal N0_29_68 : std_logic;
	signal N0_29_69 : std_logic;
	signal N0_29_70 : std_logic;
	signal N0_29_71 : std_logic;
	signal N0_29_72 : std_logic;
	signal N0_29_73 : std_logic;
	signal N0_29_74 : std_logic;
	signal N0_29_75 : std_logic;
	signal N0_29_76 : std_logic;
	signal N0_29_77 : std_logic;
	signal N0_29_78 : std_logic;
	signal N0_29_79 : std_logic;
	signal N0_29_80 : std_logic;
	signal N0_29_81 : std_logic;
	signal N0_30_30 : std_logic;
	signal N0_30_31 : std_logic;
	signal N0_30_32 : std_logic;
	signal N0_30_33 : std_logic;
	signal N0_30_34 : std_logic;
	signal N0_30_35 : std_logic;
	signal N0_30_36 : std_logic;
	signal N0_30_37 : std_logic;
	signal N0_30_38 : std_logic;
	signal N0_30_39 : std_logic;
	signal N0_30_40 : std_logic;
	signal N0_30_41 : std_logic;
	signal N0_30_42 : std_logic;
	signal N0_30_43 : std_logic;
	signal N0_30_44 : std_logic;
	signal N0_30_45 : std_logic;
	signal N0_30_46 : std_logic;
	signal N0_30_47 : std_logic;
	signal N0_30_48 : std_logic;
	signal N0_30_49 : std_logic;
	signal N0_30_50 : std_logic;
	signal N0_30_51 : std_logic;
	signal N0_30_52 : std_logic;
	signal N0_30_53 : std_logic;
	signal N0_30_54 : std_logic;
	signal N0_30_55 : std_logic;
	signal N0_30_56 : std_logic;
	signal N0_30_57 : std_logic;
	signal N0_30_58 : std_logic;
	signal N0_30_59 : std_logic;
	signal N0_30_60 : std_logic;
	signal N0_30_61 : std_logic;
	signal N0_30_62 : std_logic;
	signal N0_30_63 : std_logic;
	signal N0_30_64 : std_logic;
	signal N0_30_65 : std_logic;
	signal N0_30_66 : std_logic;
	signal N0_30_67 : std_logic;
	signal N0_30_68 : std_logic;
	signal N0_30_69 : std_logic;
	signal N0_30_70 : std_logic;
	signal N0_30_71 : std_logic;
	signal N0_30_72 : std_logic;
	signal N0_30_73 : std_logic;
	signal N0_30_74 : std_logic;
	signal N0_30_75 : std_logic;
	signal N0_30_76 : std_logic;
	signal N0_30_77 : std_logic;
	signal N0_30_78 : std_logic;
	signal N0_30_79 : std_logic;
	signal N0_30_80 : std_logic;
	signal N0_30_81 : std_logic;
	signal N0_30_82 : std_logic;
	signal N0_31_31 : std_logic;
	signal N0_31_32 : std_logic;
	signal N0_31_33 : std_logic;
	signal N0_31_34 : std_logic;
	signal N0_31_35 : std_logic;
	signal N0_31_36 : std_logic;
	signal N0_31_37 : std_logic;
	signal N0_31_38 : std_logic;
	signal N0_31_39 : std_logic;
	signal N0_31_40 : std_logic;
	signal N0_31_41 : std_logic;
	signal N0_31_42 : std_logic;
	signal N0_31_43 : std_logic;
	signal N0_31_44 : std_logic;
	signal N0_31_45 : std_logic;
	signal N0_31_46 : std_logic;
	signal N0_31_47 : std_logic;
	signal N0_31_48 : std_logic;
	signal N0_31_49 : std_logic;
	signal N0_31_50 : std_logic;
	signal N0_31_51 : std_logic;
	signal N0_31_52 : std_logic;
	signal N0_31_53 : std_logic;
	signal N0_31_54 : std_logic;
	signal N0_31_55 : std_logic;
	signal N0_31_56 : std_logic;
	signal N0_31_57 : std_logic;
	signal N0_31_58 : std_logic;
	signal N0_31_59 : std_logic;
	signal N0_31_60 : std_logic;
	signal N0_31_61 : std_logic;
	signal N0_31_62 : std_logic;
	signal N0_31_63 : std_logic;
	signal N0_31_64 : std_logic;
	signal N0_31_65 : std_logic;
	signal N0_31_66 : std_logic;
	signal N0_31_67 : std_logic;
	signal N0_31_68 : std_logic;
	signal N0_31_69 : std_logic;
	signal N0_31_70 : std_logic;
	signal N0_31_71 : std_logic;
	signal N0_31_72 : std_logic;
	signal N0_31_73 : std_logic;
	signal N0_31_74 : std_logic;
	signal N0_31_75 : std_logic;
	signal N0_31_76 : std_logic;
	signal N0_31_77 : std_logic;
	signal N0_31_78 : std_logic;
	signal N0_31_79 : std_logic;
	signal N0_31_80 : std_logic;
	signal N0_31_81 : std_logic;
	signal N0_31_82 : std_logic;
	signal N0_31_83 : std_logic;
	signal N0_32_32 : std_logic;
	signal N0_32_33 : std_logic;
	signal N0_32_34 : std_logic;
	signal N0_32_35 : std_logic;
	signal N0_32_36 : std_logic;
	signal N0_32_37 : std_logic;
	signal N0_32_38 : std_logic;
	signal N0_32_39 : std_logic;
	signal N0_32_40 : std_logic;
	signal N0_32_41 : std_logic;
	signal N0_32_42 : std_logic;
	signal N0_32_43 : std_logic;
	signal N0_32_44 : std_logic;
	signal N0_32_45 : std_logic;
	signal N0_32_46 : std_logic;
	signal N0_32_47 : std_logic;
	signal N0_32_48 : std_logic;
	signal N0_32_49 : std_logic;
	signal N0_32_50 : std_logic;
	signal N0_32_51 : std_logic;
	signal N0_32_52 : std_logic;
	signal N0_32_53 : std_logic;
	signal N0_32_54 : std_logic;
	signal N0_32_55 : std_logic;
	signal N0_32_56 : std_logic;
	signal N0_32_57 : std_logic;
	signal N0_32_58 : std_logic;
	signal N0_32_59 : std_logic;
	signal N0_32_60 : std_logic;
	signal N0_32_61 : std_logic;
	signal N0_32_62 : std_logic;
	signal N0_32_63 : std_logic;
	signal N0_32_64 : std_logic;
	signal N0_32_65 : std_logic;
	signal N0_32_66 : std_logic;
	signal N0_32_67 : std_logic;
	signal N0_32_68 : std_logic;
	signal N0_32_69 : std_logic;
	signal N0_32_70 : std_logic;
	signal N0_32_71 : std_logic;
	signal N0_32_72 : std_logic;
	signal N0_32_73 : std_logic;
	signal N0_32_74 : std_logic;
	signal N0_32_75 : std_logic;
	signal N0_32_76 : std_logic;
	signal N0_32_77 : std_logic;
	signal N0_32_78 : std_logic;
	signal N0_32_79 : std_logic;
	signal N0_32_80 : std_logic;
	signal N0_32_81 : std_logic;
	signal N0_32_82 : std_logic;
	signal N0_32_83 : std_logic;
	signal N0_32_84 : std_logic;
	signal N0_33_33 : std_logic;
	signal N0_33_34 : std_logic;
	signal N0_33_35 : std_logic;
	signal N0_33_36 : std_logic;
	signal N0_33_37 : std_logic;
	signal N0_33_38 : std_logic;
	signal N0_33_39 : std_logic;
	signal N0_33_40 : std_logic;
	signal N0_33_41 : std_logic;
	signal N0_33_42 : std_logic;
	signal N0_33_43 : std_logic;
	signal N0_33_44 : std_logic;
	signal N0_33_45 : std_logic;
	signal N0_33_46 : std_logic;
	signal N0_33_47 : std_logic;
	signal N0_33_48 : std_logic;
	signal N0_33_49 : std_logic;
	signal N0_33_50 : std_logic;
	signal N0_33_51 : std_logic;
	signal N0_33_52 : std_logic;
	signal N0_33_53 : std_logic;
	signal N0_33_54 : std_logic;
	signal N0_33_55 : std_logic;
	signal N0_33_56 : std_logic;
	signal N0_33_57 : std_logic;
	signal N0_33_58 : std_logic;
	signal N0_33_59 : std_logic;
	signal N0_33_60 : std_logic;
	signal N0_33_61 : std_logic;
	signal N0_33_62 : std_logic;
	signal N0_33_63 : std_logic;
	signal N0_33_64 : std_logic;
	signal N0_33_65 : std_logic;
	signal N0_33_66 : std_logic;
	signal N0_33_67 : std_logic;
	signal N0_33_68 : std_logic;
	signal N0_33_69 : std_logic;
	signal N0_33_70 : std_logic;
	signal N0_33_71 : std_logic;
	signal N0_33_72 : std_logic;
	signal N0_33_73 : std_logic;
	signal N0_33_74 : std_logic;
	signal N0_33_75 : std_logic;
	signal N0_33_76 : std_logic;
	signal N0_33_77 : std_logic;
	signal N0_33_78 : std_logic;
	signal N0_33_79 : std_logic;
	signal N0_33_80 : std_logic;
	signal N0_33_81 : std_logic;
	signal N0_33_82 : std_logic;
	signal N0_33_83 : std_logic;
	signal N0_33_84 : std_logic;
	signal N0_33_85 : std_logic;
	signal N0_34_34 : std_logic;
	signal N0_34_35 : std_logic;
	signal N0_34_36 : std_logic;
	signal N0_34_37 : std_logic;
	signal N0_34_38 : std_logic;
	signal N0_34_39 : std_logic;
	signal N0_34_40 : std_logic;
	signal N0_34_41 : std_logic;
	signal N0_34_42 : std_logic;
	signal N0_34_43 : std_logic;
	signal N0_34_44 : std_logic;
	signal N0_34_45 : std_logic;
	signal N0_34_46 : std_logic;
	signal N0_34_47 : std_logic;
	signal N0_34_48 : std_logic;
	signal N0_34_49 : std_logic;
	signal N0_34_50 : std_logic;
	signal N0_34_51 : std_logic;
	signal N0_34_52 : std_logic;
	signal N0_34_53 : std_logic;
	signal N0_34_54 : std_logic;
	signal N0_34_55 : std_logic;
	signal N0_34_56 : std_logic;
	signal N0_34_57 : std_logic;
	signal N0_34_58 : std_logic;
	signal N0_34_59 : std_logic;
	signal N0_34_60 : std_logic;
	signal N0_34_61 : std_logic;
	signal N0_34_62 : std_logic;
	signal N0_34_63 : std_logic;
	signal N0_34_64 : std_logic;
	signal N0_34_65 : std_logic;
	signal N0_34_66 : std_logic;
	signal N0_34_67 : std_logic;
	signal N0_34_68 : std_logic;
	signal N0_34_69 : std_logic;
	signal N0_34_70 : std_logic;
	signal N0_34_71 : std_logic;
	signal N0_34_72 : std_logic;
	signal N0_34_73 : std_logic;
	signal N0_34_74 : std_logic;
	signal N0_34_75 : std_logic;
	signal N0_34_76 : std_logic;
	signal N0_34_77 : std_logic;
	signal N0_34_78 : std_logic;
	signal N0_34_79 : std_logic;
	signal N0_34_80 : std_logic;
	signal N0_34_81 : std_logic;
	signal N0_34_82 : std_logic;
	signal N0_34_83 : std_logic;
	signal N0_34_84 : std_logic;
	signal N0_34_85 : std_logic;
	signal N0_34_86 : std_logic;
	signal N0_35_35 : std_logic;
	signal N0_35_36 : std_logic;
	signal N0_35_37 : std_logic;
	signal N0_35_38 : std_logic;
	signal N0_35_39 : std_logic;
	signal N0_35_40 : std_logic;
	signal N0_35_41 : std_logic;
	signal N0_35_42 : std_logic;
	signal N0_35_43 : std_logic;
	signal N0_35_44 : std_logic;
	signal N0_35_45 : std_logic;
	signal N0_35_46 : std_logic;
	signal N0_35_47 : std_logic;
	signal N0_35_48 : std_logic;
	signal N0_35_49 : std_logic;
	signal N0_35_50 : std_logic;
	signal N0_35_51 : std_logic;
	signal N0_35_52 : std_logic;
	signal N0_35_53 : std_logic;
	signal N0_35_54 : std_logic;
	signal N0_35_55 : std_logic;
	signal N0_35_56 : std_logic;
	signal N0_35_57 : std_logic;
	signal N0_35_58 : std_logic;
	signal N0_35_59 : std_logic;
	signal N0_35_60 : std_logic;
	signal N0_35_61 : std_logic;
	signal N0_35_62 : std_logic;
	signal N0_35_63 : std_logic;
	signal N0_35_64 : std_logic;
	signal N0_35_65 : std_logic;
	signal N0_35_66 : std_logic;
	signal N0_35_67 : std_logic;
	signal N0_35_68 : std_logic;
	signal N0_35_69 : std_logic;
	signal N0_35_70 : std_logic;
	signal N0_35_71 : std_logic;
	signal N0_35_72 : std_logic;
	signal N0_35_73 : std_logic;
	signal N0_35_74 : std_logic;
	signal N0_35_75 : std_logic;
	signal N0_35_76 : std_logic;
	signal N0_35_77 : std_logic;
	signal N0_35_78 : std_logic;
	signal N0_35_79 : std_logic;
	signal N0_35_80 : std_logic;
	signal N0_35_81 : std_logic;
	signal N0_35_82 : std_logic;
	signal N0_35_83 : std_logic;
	signal N0_35_84 : std_logic;
	signal N0_35_85 : std_logic;
	signal N0_35_86 : std_logic;
	signal N0_35_87 : std_logic;
	signal N0_36_36 : std_logic;
	signal N0_36_37 : std_logic;
	signal N0_36_38 : std_logic;
	signal N0_36_39 : std_logic;
	signal N0_36_40 : std_logic;
	signal N0_36_41 : std_logic;
	signal N0_36_42 : std_logic;
	signal N0_36_43 : std_logic;
	signal N0_36_44 : std_logic;
	signal N0_36_45 : std_logic;
	signal N0_36_46 : std_logic;
	signal N0_36_47 : std_logic;
	signal N0_36_48 : std_logic;
	signal N0_36_49 : std_logic;
	signal N0_36_50 : std_logic;
	signal N0_36_51 : std_logic;
	signal N0_36_52 : std_logic;
	signal N0_36_53 : std_logic;
	signal N0_36_54 : std_logic;
	signal N0_36_55 : std_logic;
	signal N0_36_56 : std_logic;
	signal N0_36_57 : std_logic;
	signal N0_36_58 : std_logic;
	signal N0_36_59 : std_logic;
	signal N0_36_60 : std_logic;
	signal N0_36_61 : std_logic;
	signal N0_36_62 : std_logic;
	signal N0_36_63 : std_logic;
	signal N0_36_64 : std_logic;
	signal N0_36_65 : std_logic;
	signal N0_36_66 : std_logic;
	signal N0_36_67 : std_logic;
	signal N0_36_68 : std_logic;
	signal N0_36_69 : std_logic;
	signal N0_36_70 : std_logic;
	signal N0_36_71 : std_logic;
	signal N0_36_72 : std_logic;
	signal N0_36_73 : std_logic;
	signal N0_36_74 : std_logic;
	signal N0_36_75 : std_logic;
	signal N0_36_76 : std_logic;
	signal N0_36_77 : std_logic;
	signal N0_36_78 : std_logic;
	signal N0_36_79 : std_logic;
	signal N0_36_80 : std_logic;
	signal N0_36_81 : std_logic;
	signal N0_36_82 : std_logic;
	signal N0_36_83 : std_logic;
	signal N0_36_84 : std_logic;
	signal N0_36_85 : std_logic;
	signal N0_36_86 : std_logic;
	signal N0_36_87 : std_logic;
	signal N0_36_88 : std_logic;
	signal N0_37_37 : std_logic;
	signal N0_37_38 : std_logic;
	signal N0_37_39 : std_logic;
	signal N0_37_40 : std_logic;
	signal N0_37_41 : std_logic;
	signal N0_37_42 : std_logic;
	signal N0_37_43 : std_logic;
	signal N0_37_44 : std_logic;
	signal N0_37_45 : std_logic;
	signal N0_37_46 : std_logic;
	signal N0_37_47 : std_logic;
	signal N0_37_48 : std_logic;
	signal N0_37_49 : std_logic;
	signal N0_37_50 : std_logic;
	signal N0_37_51 : std_logic;
	signal N0_37_52 : std_logic;
	signal N0_37_53 : std_logic;
	signal N0_37_54 : std_logic;
	signal N0_37_55 : std_logic;
	signal N0_37_56 : std_logic;
	signal N0_37_57 : std_logic;
	signal N0_37_58 : std_logic;
	signal N0_37_59 : std_logic;
	signal N0_37_60 : std_logic;
	signal N0_37_61 : std_logic;
	signal N0_37_62 : std_logic;
	signal N0_37_63 : std_logic;
	signal N0_37_64 : std_logic;
	signal N0_37_65 : std_logic;
	signal N0_37_66 : std_logic;
	signal N0_37_67 : std_logic;
	signal N0_37_68 : std_logic;
	signal N0_37_69 : std_logic;
	signal N0_37_70 : std_logic;
	signal N0_37_71 : std_logic;
	signal N0_37_72 : std_logic;
	signal N0_37_73 : std_logic;
	signal N0_37_74 : std_logic;
	signal N0_37_75 : std_logic;
	signal N0_37_76 : std_logic;
	signal N0_37_77 : std_logic;
	signal N0_37_78 : std_logic;
	signal N0_37_79 : std_logic;
	signal N0_37_80 : std_logic;
	signal N0_37_81 : std_logic;
	signal N0_37_82 : std_logic;
	signal N0_37_83 : std_logic;
	signal N0_37_84 : std_logic;
	signal N0_37_85 : std_logic;
	signal N0_37_86 : std_logic;
	signal N0_37_87 : std_logic;
	signal N0_37_88 : std_logic;
	signal N0_37_89 : std_logic;
	signal N0_38_38 : std_logic;
	signal N0_38_39 : std_logic;
	signal N0_38_40 : std_logic;
	signal N0_38_41 : std_logic;
	signal N0_38_42 : std_logic;
	signal N0_38_43 : std_logic;
	signal N0_38_44 : std_logic;
	signal N0_38_45 : std_logic;
	signal N0_38_46 : std_logic;
	signal N0_38_47 : std_logic;
	signal N0_38_48 : std_logic;
	signal N0_38_49 : std_logic;
	signal N0_38_50 : std_logic;
	signal N0_38_51 : std_logic;
	signal N0_38_52 : std_logic;
	signal N0_38_53 : std_logic;
	signal N0_38_54 : std_logic;
	signal N0_38_55 : std_logic;
	signal N0_38_56 : std_logic;
	signal N0_38_57 : std_logic;
	signal N0_38_58 : std_logic;
	signal N0_38_59 : std_logic;
	signal N0_38_60 : std_logic;
	signal N0_38_61 : std_logic;
	signal N0_38_62 : std_logic;
	signal N0_38_63 : std_logic;
	signal N0_38_64 : std_logic;
	signal N0_38_65 : std_logic;
	signal N0_38_66 : std_logic;
	signal N0_38_67 : std_logic;
	signal N0_38_68 : std_logic;
	signal N0_38_69 : std_logic;
	signal N0_38_70 : std_logic;
	signal N0_38_71 : std_logic;
	signal N0_38_72 : std_logic;
	signal N0_38_73 : std_logic;
	signal N0_38_74 : std_logic;
	signal N0_38_75 : std_logic;
	signal N0_38_76 : std_logic;
	signal N0_38_77 : std_logic;
	signal N0_38_78 : std_logic;
	signal N0_38_79 : std_logic;
	signal N0_38_80 : std_logic;
	signal N0_38_81 : std_logic;
	signal N0_38_82 : std_logic;
	signal N0_38_83 : std_logic;
	signal N0_38_84 : std_logic;
	signal N0_38_85 : std_logic;
	signal N0_38_86 : std_logic;
	signal N0_38_87 : std_logic;
	signal N0_38_88 : std_logic;
	signal N0_38_89 : std_logic;
	signal N0_38_90 : std_logic;
	signal N0_39_39 : std_logic;
	signal N0_39_40 : std_logic;
	signal N0_39_41 : std_logic;
	signal N0_39_42 : std_logic;
	signal N0_39_43 : std_logic;
	signal N0_39_44 : std_logic;
	signal N0_39_45 : std_logic;
	signal N0_39_46 : std_logic;
	signal N0_39_47 : std_logic;
	signal N0_39_48 : std_logic;
	signal N0_39_49 : std_logic;
	signal N0_39_50 : std_logic;
	signal N0_39_51 : std_logic;
	signal N0_39_52 : std_logic;
	signal N0_39_53 : std_logic;
	signal N0_39_54 : std_logic;
	signal N0_39_55 : std_logic;
	signal N0_39_56 : std_logic;
	signal N0_39_57 : std_logic;
	signal N0_39_58 : std_logic;
	signal N0_39_59 : std_logic;
	signal N0_39_60 : std_logic;
	signal N0_39_61 : std_logic;
	signal N0_39_62 : std_logic;
	signal N0_39_63 : std_logic;
	signal N0_39_64 : std_logic;
	signal N0_39_65 : std_logic;
	signal N0_39_66 : std_logic;
	signal N0_39_67 : std_logic;
	signal N0_39_68 : std_logic;
	signal N0_39_69 : std_logic;
	signal N0_39_70 : std_logic;
	signal N0_39_71 : std_logic;
	signal N0_39_72 : std_logic;
	signal N0_39_73 : std_logic;
	signal N0_39_74 : std_logic;
	signal N0_39_75 : std_logic;
	signal N0_39_76 : std_logic;
	signal N0_39_77 : std_logic;
	signal N0_39_78 : std_logic;
	signal N0_39_79 : std_logic;
	signal N0_39_80 : std_logic;
	signal N0_39_81 : std_logic;
	signal N0_39_82 : std_logic;
	signal N0_39_83 : std_logic;
	signal N0_39_84 : std_logic;
	signal N0_39_85 : std_logic;
	signal N0_39_86 : std_logic;
	signal N0_39_87 : std_logic;
	signal N0_39_88 : std_logic;
	signal N0_39_89 : std_logic;
	signal N0_39_90 : std_logic;
	signal N0_39_91 : std_logic;
	signal N0_40_40 : std_logic;
	signal N0_40_41 : std_logic;
	signal N0_40_42 : std_logic;
	signal N0_40_43 : std_logic;
	signal N0_40_44 : std_logic;
	signal N0_40_45 : std_logic;
	signal N0_40_46 : std_logic;
	signal N0_40_47 : std_logic;
	signal N0_40_48 : std_logic;
	signal N0_40_49 : std_logic;
	signal N0_40_50 : std_logic;
	signal N0_40_51 : std_logic;
	signal N0_40_52 : std_logic;
	signal N0_40_53 : std_logic;
	signal N0_40_54 : std_logic;
	signal N0_40_55 : std_logic;
	signal N0_40_56 : std_logic;
	signal N0_40_57 : std_logic;
	signal N0_40_58 : std_logic;
	signal N0_40_59 : std_logic;
	signal N0_40_60 : std_logic;
	signal N0_40_61 : std_logic;
	signal N0_40_62 : std_logic;
	signal N0_40_63 : std_logic;
	signal N0_40_64 : std_logic;
	signal N0_40_65 : std_logic;
	signal N0_40_66 : std_logic;
	signal N0_40_67 : std_logic;
	signal N0_40_68 : std_logic;
	signal N0_40_69 : std_logic;
	signal N0_40_70 : std_logic;
	signal N0_40_71 : std_logic;
	signal N0_40_72 : std_logic;
	signal N0_40_73 : std_logic;
	signal N0_40_74 : std_logic;
	signal N0_40_75 : std_logic;
	signal N0_40_76 : std_logic;
	signal N0_40_77 : std_logic;
	signal N0_40_78 : std_logic;
	signal N0_40_79 : std_logic;
	signal N0_40_80 : std_logic;
	signal N0_40_81 : std_logic;
	signal N0_40_82 : std_logic;
	signal N0_40_83 : std_logic;
	signal N0_40_84 : std_logic;
	signal N0_40_85 : std_logic;
	signal N0_40_86 : std_logic;
	signal N0_40_87 : std_logic;
	signal N0_40_88 : std_logic;
	signal N0_40_89 : std_logic;
	signal N0_40_90 : std_logic;
	signal N0_40_91 : std_logic;
	signal N0_40_92 : std_logic;
	signal N0_41_41 : std_logic;
	signal N0_41_42 : std_logic;
	signal N0_41_43 : std_logic;
	signal N0_41_44 : std_logic;
	signal N0_41_45 : std_logic;
	signal N0_41_46 : std_logic;
	signal N0_41_47 : std_logic;
	signal N0_41_48 : std_logic;
	signal N0_41_49 : std_logic;
	signal N0_41_50 : std_logic;
	signal N0_41_51 : std_logic;
	signal N0_41_52 : std_logic;
	signal N0_41_53 : std_logic;
	signal N0_41_54 : std_logic;
	signal N0_41_55 : std_logic;
	signal N0_41_56 : std_logic;
	signal N0_41_57 : std_logic;
	signal N0_41_58 : std_logic;
	signal N0_41_59 : std_logic;
	signal N0_41_60 : std_logic;
	signal N0_41_61 : std_logic;
	signal N0_41_62 : std_logic;
	signal N0_41_63 : std_logic;
	signal N0_41_64 : std_logic;
	signal N0_41_65 : std_logic;
	signal N0_41_66 : std_logic;
	signal N0_41_67 : std_logic;
	signal N0_41_68 : std_logic;
	signal N0_41_69 : std_logic;
	signal N0_41_70 : std_logic;
	signal N0_41_71 : std_logic;
	signal N0_41_72 : std_logic;
	signal N0_41_73 : std_logic;
	signal N0_41_74 : std_logic;
	signal N0_41_75 : std_logic;
	signal N0_41_76 : std_logic;
	signal N0_41_77 : std_logic;
	signal N0_41_78 : std_logic;
	signal N0_41_79 : std_logic;
	signal N0_41_80 : std_logic;
	signal N0_41_81 : std_logic;
	signal N0_41_82 : std_logic;
	signal N0_41_83 : std_logic;
	signal N0_41_84 : std_logic;
	signal N0_41_85 : std_logic;
	signal N0_41_86 : std_logic;
	signal N0_41_87 : std_logic;
	signal N0_41_88 : std_logic;
	signal N0_41_89 : std_logic;
	signal N0_41_90 : std_logic;
	signal N0_41_91 : std_logic;
	signal N0_41_92 : std_logic;
	signal N0_41_93 : std_logic;
	signal N0_42_42 : std_logic;
	signal N0_42_43 : std_logic;
	signal N0_42_44 : std_logic;
	signal N0_42_45 : std_logic;
	signal N0_42_46 : std_logic;
	signal N0_42_47 : std_logic;
	signal N0_42_48 : std_logic;
	signal N0_42_49 : std_logic;
	signal N0_42_50 : std_logic;
	signal N0_42_51 : std_logic;
	signal N0_42_52 : std_logic;
	signal N0_42_53 : std_logic;
	signal N0_42_54 : std_logic;
	signal N0_42_55 : std_logic;
	signal N0_42_56 : std_logic;
	signal N0_42_57 : std_logic;
	signal N0_42_58 : std_logic;
	signal N0_42_59 : std_logic;
	signal N0_42_60 : std_logic;
	signal N0_42_61 : std_logic;
	signal N0_42_62 : std_logic;
	signal N0_42_63 : std_logic;
	signal N0_42_64 : std_logic;
	signal N0_42_65 : std_logic;
	signal N0_42_66 : std_logic;
	signal N0_42_67 : std_logic;
	signal N0_42_68 : std_logic;
	signal N0_42_69 : std_logic;
	signal N0_42_70 : std_logic;
	signal N0_42_71 : std_logic;
	signal N0_42_72 : std_logic;
	signal N0_42_73 : std_logic;
	signal N0_42_74 : std_logic;
	signal N0_42_75 : std_logic;
	signal N0_42_76 : std_logic;
	signal N0_42_77 : std_logic;
	signal N0_42_78 : std_logic;
	signal N0_42_79 : std_logic;
	signal N0_42_80 : std_logic;
	signal N0_42_81 : std_logic;
	signal N0_42_82 : std_logic;
	signal N0_42_83 : std_logic;
	signal N0_42_84 : std_logic;
	signal N0_42_85 : std_logic;
	signal N0_42_86 : std_logic;
	signal N0_42_87 : std_logic;
	signal N0_42_88 : std_logic;
	signal N0_42_89 : std_logic;
	signal N0_42_90 : std_logic;
	signal N0_42_91 : std_logic;
	signal N0_42_92 : std_logic;
	signal N0_42_93 : std_logic;
	signal N0_42_94 : std_logic;
	signal N0_43_43 : std_logic;
	signal N0_43_44 : std_logic;
	signal N0_43_45 : std_logic;
	signal N0_43_46 : std_logic;
	signal N0_43_47 : std_logic;
	signal N0_43_48 : std_logic;
	signal N0_43_49 : std_logic;
	signal N0_43_50 : std_logic;
	signal N0_43_51 : std_logic;
	signal N0_43_52 : std_logic;
	signal N0_43_53 : std_logic;
	signal N0_43_54 : std_logic;
	signal N0_43_55 : std_logic;
	signal N0_43_56 : std_logic;
	signal N0_43_57 : std_logic;
	signal N0_43_58 : std_logic;
	signal N0_43_59 : std_logic;
	signal N0_43_60 : std_logic;
	signal N0_43_61 : std_logic;
	signal N0_43_62 : std_logic;
	signal N0_43_63 : std_logic;
	signal N0_43_64 : std_logic;
	signal N0_43_65 : std_logic;
	signal N0_43_66 : std_logic;
	signal N0_43_67 : std_logic;
	signal N0_43_68 : std_logic;
	signal N0_43_69 : std_logic;
	signal N0_43_70 : std_logic;
	signal N0_43_71 : std_logic;
	signal N0_43_72 : std_logic;
	signal N0_43_73 : std_logic;
	signal N0_43_74 : std_logic;
	signal N0_43_75 : std_logic;
	signal N0_43_76 : std_logic;
	signal N0_43_77 : std_logic;
	signal N0_43_78 : std_logic;
	signal N0_43_79 : std_logic;
	signal N0_43_80 : std_logic;
	signal N0_43_81 : std_logic;
	signal N0_43_82 : std_logic;
	signal N0_43_83 : std_logic;
	signal N0_43_84 : std_logic;
	signal N0_43_85 : std_logic;
	signal N0_43_86 : std_logic;
	signal N0_43_87 : std_logic;
	signal N0_43_88 : std_logic;
	signal N0_43_89 : std_logic;
	signal N0_43_90 : std_logic;
	signal N0_43_91 : std_logic;
	signal N0_43_92 : std_logic;
	signal N0_43_93 : std_logic;
	signal N0_43_94 : std_logic;
	signal N0_43_95 : std_logic;
	signal N0_44_44 : std_logic;
	signal N0_44_45 : std_logic;
	signal N0_44_46 : std_logic;
	signal N0_44_47 : std_logic;
	signal N0_44_48 : std_logic;
	signal N0_44_49 : std_logic;
	signal N0_44_50 : std_logic;
	signal N0_44_51 : std_logic;
	signal N0_44_52 : std_logic;
	signal N0_44_53 : std_logic;
	signal N0_44_54 : std_logic;
	signal N0_44_55 : std_logic;
	signal N0_44_56 : std_logic;
	signal N0_44_57 : std_logic;
	signal N0_44_58 : std_logic;
	signal N0_44_59 : std_logic;
	signal N0_44_60 : std_logic;
	signal N0_44_61 : std_logic;
	signal N0_44_62 : std_logic;
	signal N0_44_63 : std_logic;
	signal N0_44_64 : std_logic;
	signal N0_44_65 : std_logic;
	signal N0_44_66 : std_logic;
	signal N0_44_67 : std_logic;
	signal N0_44_68 : std_logic;
	signal N0_44_69 : std_logic;
	signal N0_44_70 : std_logic;
	signal N0_44_71 : std_logic;
	signal N0_44_72 : std_logic;
	signal N0_44_73 : std_logic;
	signal N0_44_74 : std_logic;
	signal N0_44_75 : std_logic;
	signal N0_44_76 : std_logic;
	signal N0_44_77 : std_logic;
	signal N0_44_78 : std_logic;
	signal N0_44_79 : std_logic;
	signal N0_44_80 : std_logic;
	signal N0_44_81 : std_logic;
	signal N0_44_82 : std_logic;
	signal N0_44_83 : std_logic;
	signal N0_44_84 : std_logic;
	signal N0_44_85 : std_logic;
	signal N0_44_86 : std_logic;
	signal N0_44_87 : std_logic;
	signal N0_44_88 : std_logic;
	signal N0_44_89 : std_logic;
	signal N0_44_90 : std_logic;
	signal N0_44_91 : std_logic;
	signal N0_44_92 : std_logic;
	signal N0_44_93 : std_logic;
	signal N0_44_94 : std_logic;
	signal N0_44_95 : std_logic;
	signal N0_44_96 : std_logic;
	signal N0_45_45 : std_logic;
	signal N0_45_46 : std_logic;
	signal N0_45_47 : std_logic;
	signal N0_45_48 : std_logic;
	signal N0_45_49 : std_logic;
	signal N0_45_50 : std_logic;
	signal N0_45_51 : std_logic;
	signal N0_45_52 : std_logic;
	signal N0_45_53 : std_logic;
	signal N0_45_54 : std_logic;
	signal N0_45_55 : std_logic;
	signal N0_45_56 : std_logic;
	signal N0_45_57 : std_logic;
	signal N0_45_58 : std_logic;
	signal N0_45_59 : std_logic;
	signal N0_45_60 : std_logic;
	signal N0_45_61 : std_logic;
	signal N0_45_62 : std_logic;
	signal N0_45_63 : std_logic;
	signal N0_45_64 : std_logic;
	signal N0_45_65 : std_logic;
	signal N0_45_66 : std_logic;
	signal N0_45_67 : std_logic;
	signal N0_45_68 : std_logic;
	signal N0_45_69 : std_logic;
	signal N0_45_70 : std_logic;
	signal N0_45_71 : std_logic;
	signal N0_45_72 : std_logic;
	signal N0_45_73 : std_logic;
	signal N0_45_74 : std_logic;
	signal N0_45_75 : std_logic;
	signal N0_45_76 : std_logic;
	signal N0_45_77 : std_logic;
	signal N0_45_78 : std_logic;
	signal N0_45_79 : std_logic;
	signal N0_45_80 : std_logic;
	signal N0_45_81 : std_logic;
	signal N0_45_82 : std_logic;
	signal N0_45_83 : std_logic;
	signal N0_45_84 : std_logic;
	signal N0_45_85 : std_logic;
	signal N0_45_86 : std_logic;
	signal N0_45_87 : std_logic;
	signal N0_45_88 : std_logic;
	signal N0_45_89 : std_logic;
	signal N0_45_90 : std_logic;
	signal N0_45_91 : std_logic;
	signal N0_45_92 : std_logic;
	signal N0_45_93 : std_logic;
	signal N0_45_94 : std_logic;
	signal N0_45_95 : std_logic;
	signal N0_45_96 : std_logic;
	signal N0_45_97 : std_logic;
	signal N0_46_46 : std_logic;
	signal N0_46_47 : std_logic;
	signal N0_46_48 : std_logic;
	signal N0_46_49 : std_logic;
	signal N0_46_50 : std_logic;
	signal N0_46_51 : std_logic;
	signal N0_46_52 : std_logic;
	signal N0_46_53 : std_logic;
	signal N0_46_54 : std_logic;
	signal N0_46_55 : std_logic;
	signal N0_46_56 : std_logic;
	signal N0_46_57 : std_logic;
	signal N0_46_58 : std_logic;
	signal N0_46_59 : std_logic;
	signal N0_46_60 : std_logic;
	signal N0_46_61 : std_logic;
	signal N0_46_62 : std_logic;
	signal N0_46_63 : std_logic;
	signal N0_46_64 : std_logic;
	signal N0_46_65 : std_logic;
	signal N0_46_66 : std_logic;
	signal N0_46_67 : std_logic;
	signal N0_46_68 : std_logic;
	signal N0_46_69 : std_logic;
	signal N0_46_70 : std_logic;
	signal N0_46_71 : std_logic;
	signal N0_46_72 : std_logic;
	signal N0_46_73 : std_logic;
	signal N0_46_74 : std_logic;
	signal N0_46_75 : std_logic;
	signal N0_46_76 : std_logic;
	signal N0_46_77 : std_logic;
	signal N0_46_78 : std_logic;
	signal N0_46_79 : std_logic;
	signal N0_46_80 : std_logic;
	signal N0_46_81 : std_logic;
	signal N0_46_82 : std_logic;
	signal N0_46_83 : std_logic;
	signal N0_46_84 : std_logic;
	signal N0_46_85 : std_logic;
	signal N0_46_86 : std_logic;
	signal N0_46_87 : std_logic;
	signal N0_46_88 : std_logic;
	signal N0_46_89 : std_logic;
	signal N0_46_90 : std_logic;
	signal N0_46_91 : std_logic;
	signal N0_46_92 : std_logic;
	signal N0_46_93 : std_logic;
	signal N0_46_94 : std_logic;
	signal N0_46_95 : std_logic;
	signal N0_46_96 : std_logic;
	signal N0_46_97 : std_logic;
	signal N0_46_98 : std_logic;
	signal N0_47_47 : std_logic;
	signal N0_47_48 : std_logic;
	signal N0_47_49 : std_logic;
	signal N0_47_50 : std_logic;
	signal N0_47_51 : std_logic;
	signal N0_47_52 : std_logic;
	signal N0_47_53 : std_logic;
	signal N0_47_54 : std_logic;
	signal N0_47_55 : std_logic;
	signal N0_47_56 : std_logic;
	signal N0_47_57 : std_logic;
	signal N0_47_58 : std_logic;
	signal N0_47_59 : std_logic;
	signal N0_47_60 : std_logic;
	signal N0_47_61 : std_logic;
	signal N0_47_62 : std_logic;
	signal N0_47_63 : std_logic;
	signal N0_47_64 : std_logic;
	signal N0_47_65 : std_logic;
	signal N0_47_66 : std_logic;
	signal N0_47_67 : std_logic;
	signal N0_47_68 : std_logic;
	signal N0_47_69 : std_logic;
	signal N0_47_70 : std_logic;
	signal N0_47_71 : std_logic;
	signal N0_47_72 : std_logic;
	signal N0_47_73 : std_logic;
	signal N0_47_74 : std_logic;
	signal N0_47_75 : std_logic;
	signal N0_47_76 : std_logic;
	signal N0_47_77 : std_logic;
	signal N0_47_78 : std_logic;
	signal N0_47_79 : std_logic;
	signal N0_47_80 : std_logic;
	signal N0_47_81 : std_logic;
	signal N0_47_82 : std_logic;
	signal N0_47_83 : std_logic;
	signal N0_47_84 : std_logic;
	signal N0_47_85 : std_logic;
	signal N0_47_86 : std_logic;
	signal N0_47_87 : std_logic;
	signal N0_47_88 : std_logic;
	signal N0_47_89 : std_logic;
	signal N0_47_90 : std_logic;
	signal N0_47_91 : std_logic;
	signal N0_47_92 : std_logic;
	signal N0_47_93 : std_logic;
	signal N0_47_94 : std_logic;
	signal N0_47_95 : std_logic;
	signal N0_47_96 : std_logic;
	signal N0_47_97 : std_logic;
	signal N0_47_98 : std_logic;
	signal N0_47_99 : std_logic;
	signal N0_48_48 : std_logic;
	signal N0_48_49 : std_logic;
	signal N0_48_50 : std_logic;
	signal N0_48_51 : std_logic;
	signal N0_48_52 : std_logic;
	signal N0_48_53 : std_logic;
	signal N0_48_54 : std_logic;
	signal N0_48_55 : std_logic;
	signal N0_48_56 : std_logic;
	signal N0_48_57 : std_logic;
	signal N0_48_58 : std_logic;
	signal N0_48_59 : std_logic;
	signal N0_48_60 : std_logic;
	signal N0_48_61 : std_logic;
	signal N0_48_62 : std_logic;
	signal N0_48_63 : std_logic;
	signal N0_48_64 : std_logic;
	signal N0_48_65 : std_logic;
	signal N0_48_66 : std_logic;
	signal N0_48_67 : std_logic;
	signal N0_48_68 : std_logic;
	signal N0_48_69 : std_logic;
	signal N0_48_70 : std_logic;
	signal N0_48_71 : std_logic;
	signal N0_48_72 : std_logic;
	signal N0_48_73 : std_logic;
	signal N0_48_74 : std_logic;
	signal N0_48_75 : std_logic;
	signal N0_48_76 : std_logic;
	signal N0_48_77 : std_logic;
	signal N0_48_78 : std_logic;
	signal N0_48_79 : std_logic;
	signal N0_48_80 : std_logic;
	signal N0_48_81 : std_logic;
	signal N0_48_82 : std_logic;
	signal N0_48_83 : std_logic;
	signal N0_48_84 : std_logic;
	signal N0_48_85 : std_logic;
	signal N0_48_86 : std_logic;
	signal N0_48_87 : std_logic;
	signal N0_48_88 : std_logic;
	signal N0_48_89 : std_logic;
	signal N0_48_90 : std_logic;
	signal N0_48_91 : std_logic;
	signal N0_48_92 : std_logic;
	signal N0_48_93 : std_logic;
	signal N0_48_94 : std_logic;
	signal N0_48_95 : std_logic;
	signal N0_48_96 : std_logic;
	signal N0_48_97 : std_logic;
	signal N0_48_98 : std_logic;
	signal N0_48_99 : std_logic;
	signal N0_48_100 : std_logic;
	signal N0_49_49 : std_logic;
	signal N0_49_50 : std_logic;
	signal N0_49_51 : std_logic;
	signal N0_49_52 : std_logic;
	signal N0_49_53 : std_logic;
	signal N0_49_54 : std_logic;
	signal N0_49_55 : std_logic;
	signal N0_49_56 : std_logic;
	signal N0_49_57 : std_logic;
	signal N0_49_58 : std_logic;
	signal N0_49_59 : std_logic;
	signal N0_49_60 : std_logic;
	signal N0_49_61 : std_logic;
	signal N0_49_62 : std_logic;
	signal N0_49_63 : std_logic;
	signal N0_49_64 : std_logic;
	signal N0_49_65 : std_logic;
	signal N0_49_66 : std_logic;
	signal N0_49_67 : std_logic;
	signal N0_49_68 : std_logic;
	signal N0_49_69 : std_logic;
	signal N0_49_70 : std_logic;
	signal N0_49_71 : std_logic;
	signal N0_49_72 : std_logic;
	signal N0_49_73 : std_logic;
	signal N0_49_74 : std_logic;
	signal N0_49_75 : std_logic;
	signal N0_49_76 : std_logic;
	signal N0_49_77 : std_logic;
	signal N0_49_78 : std_logic;
	signal N0_49_79 : std_logic;
	signal N0_49_80 : std_logic;
	signal N0_49_81 : std_logic;
	signal N0_49_82 : std_logic;
	signal N0_49_83 : std_logic;
	signal N0_49_84 : std_logic;
	signal N0_49_85 : std_logic;
	signal N0_49_86 : std_logic;
	signal N0_49_87 : std_logic;
	signal N0_49_88 : std_logic;
	signal N0_49_89 : std_logic;
	signal N0_49_90 : std_logic;
	signal N0_49_91 : std_logic;
	signal N0_49_92 : std_logic;
	signal N0_49_93 : std_logic;
	signal N0_49_94 : std_logic;
	signal N0_49_95 : std_logic;
	signal N0_49_96 : std_logic;
	signal N0_49_97 : std_logic;
	signal N0_49_98 : std_logic;
	signal N0_49_99 : std_logic;
	signal N0_49_100 : std_logic;
	signal N0_49_101 : std_logic;
	signal N0_50_50 : std_logic;
	signal N0_50_51 : std_logic;
	signal N0_50_52 : std_logic;
	signal N0_50_53 : std_logic;
	signal N0_50_54 : std_logic;
	signal N0_50_55 : std_logic;
	signal N0_50_56 : std_logic;
	signal N0_50_57 : std_logic;
	signal N0_50_58 : std_logic;
	signal N0_50_59 : std_logic;
	signal N0_50_60 : std_logic;
	signal N0_50_61 : std_logic;
	signal N0_50_62 : std_logic;
	signal N0_50_63 : std_logic;
	signal N0_50_64 : std_logic;
	signal N0_50_65 : std_logic;
	signal N0_50_66 : std_logic;
	signal N0_50_67 : std_logic;
	signal N0_50_68 : std_logic;
	signal N0_50_69 : std_logic;
	signal N0_50_70 : std_logic;
	signal N0_50_71 : std_logic;
	signal N0_50_72 : std_logic;
	signal N0_50_73 : std_logic;
	signal N0_50_74 : std_logic;
	signal N0_50_75 : std_logic;
	signal N0_50_76 : std_logic;
	signal N0_50_77 : std_logic;
	signal N0_50_78 : std_logic;
	signal N0_50_79 : std_logic;
	signal N0_50_80 : std_logic;
	signal N0_50_81 : std_logic;
	signal N0_50_82 : std_logic;
	signal N0_50_83 : std_logic;
	signal N0_50_84 : std_logic;
	signal N0_50_85 : std_logic;
	signal N0_50_86 : std_logic;
	signal N0_50_87 : std_logic;
	signal N0_50_88 : std_logic;
	signal N0_50_89 : std_logic;
	signal N0_50_90 : std_logic;
	signal N0_50_91 : std_logic;
	signal N0_50_92 : std_logic;
	signal N0_50_93 : std_logic;
	signal N0_50_94 : std_logic;
	signal N0_50_95 : std_logic;
	signal N0_50_96 : std_logic;
	signal N0_50_97 : std_logic;
	signal N0_50_98 : std_logic;
	signal N0_50_99 : std_logic;
	signal N0_50_100 : std_logic;
	signal N0_50_101 : std_logic;
	signal N0_50_102 : std_logic;
	signal N0_51_51 : std_logic;
	signal N0_51_52 : std_logic;
	signal N0_51_53 : std_logic;
	signal N0_51_54 : std_logic;
	signal N0_51_55 : std_logic;
	signal N0_51_56 : std_logic;
	signal N0_51_57 : std_logic;
	signal N0_51_58 : std_logic;
	signal N0_51_59 : std_logic;
	signal N0_51_60 : std_logic;
	signal N0_51_61 : std_logic;
	signal N0_51_62 : std_logic;
	signal N0_51_63 : std_logic;
	signal N0_51_64 : std_logic;
	signal N0_51_65 : std_logic;
	signal N0_51_66 : std_logic;
	signal N0_51_67 : std_logic;
	signal N0_51_68 : std_logic;
	signal N0_51_69 : std_logic;
	signal N0_51_70 : std_logic;
	signal N0_51_71 : std_logic;
	signal N0_51_72 : std_logic;
	signal N0_51_73 : std_logic;
	signal N0_51_74 : std_logic;
	signal N0_51_75 : std_logic;
	signal N0_51_76 : std_logic;
	signal N0_51_77 : std_logic;
	signal N0_51_78 : std_logic;
	signal N0_51_79 : std_logic;
	signal N0_51_80 : std_logic;
	signal N0_51_81 : std_logic;
	signal N0_51_82 : std_logic;
	signal N0_51_83 : std_logic;
	signal N0_51_84 : std_logic;
	signal N0_51_85 : std_logic;
	signal N0_51_86 : std_logic;
	signal N0_51_87 : std_logic;
	signal N0_51_88 : std_logic;
	signal N0_51_89 : std_logic;
	signal N0_51_90 : std_logic;
	signal N0_51_91 : std_logic;
	signal N0_51_92 : std_logic;
	signal N0_51_93 : std_logic;
	signal N0_51_94 : std_logic;
	signal N0_51_95 : std_logic;
	signal N0_51_96 : std_logic;
	signal N0_51_97 : std_logic;
	signal N0_51_98 : std_logic;
	signal N0_51_99 : std_logic;
	signal N0_51_100 : std_logic;
	signal N0_51_101 : std_logic;
	signal N0_51_102 : std_logic;
	signal N0_51_103 : std_logic;
	signal N0_52_52 : std_logic;
	signal N0_52_53 : std_logic;
	signal N0_52_54 : std_logic;
	signal N0_52_55 : std_logic;
	signal N0_52_56 : std_logic;
	signal N0_52_57 : std_logic;
	signal N0_52_58 : std_logic;
	signal N0_52_59 : std_logic;
	signal N0_52_60 : std_logic;
	signal N0_52_61 : std_logic;
	signal N0_52_62 : std_logic;
	signal N0_52_63 : std_logic;
	signal N0_52_64 : std_logic;
	signal N0_52_65 : std_logic;
	signal N0_52_66 : std_logic;
	signal N0_52_67 : std_logic;
	signal N0_52_68 : std_logic;
	signal N0_52_69 : std_logic;
	signal N0_52_70 : std_logic;
	signal N0_52_71 : std_logic;
	signal N0_52_72 : std_logic;
	signal N0_52_73 : std_logic;
	signal N0_52_74 : std_logic;
	signal N0_52_75 : std_logic;
	signal N0_52_76 : std_logic;
	signal N0_52_77 : std_logic;
	signal N0_52_78 : std_logic;
	signal N0_52_79 : std_logic;
	signal N0_52_80 : std_logic;
	signal N0_52_81 : std_logic;
	signal N0_52_82 : std_logic;
	signal N0_52_83 : std_logic;
	signal N0_52_84 : std_logic;
	signal N0_52_85 : std_logic;
	signal N0_52_86 : std_logic;
	signal N0_52_87 : std_logic;
	signal N0_52_88 : std_logic;
	signal N0_52_89 : std_logic;
	signal N0_52_90 : std_logic;
	signal N0_52_91 : std_logic;
	signal N0_52_92 : std_logic;
	signal N0_52_93 : std_logic;
	signal N0_52_94 : std_logic;
	signal N0_52_95 : std_logic;
	signal N0_52_96 : std_logic;
	signal N0_52_97 : std_logic;
	signal N0_52_98 : std_logic;
	signal N0_52_99 : std_logic;
	signal N0_52_100 : std_logic;
	signal N0_52_101 : std_logic;
	signal N0_52_102 : std_logic;
	signal N0_52_103 : std_logic;
	signal N0_52_104 : std_logic;
	signal N2_0_36 : std_logic;
	signal N2_1_37 : std_logic;
	signal N2_0_37 : std_logic;
	signal N2_1_38 : std_logic;
	signal N2_2_37 : std_logic;
	signal N2_3_38 : std_logic;
	signal N2_0_38 : std_logic;
	signal N2_1_39 : std_logic;
	signal N2_2_38 : std_logic;
	signal N2_3_39 : std_logic;
	signal N2_4_38 : std_logic;
	signal N2_5_39 : std_logic;
	signal N2_0_39 : std_logic;
	signal N2_1_40 : std_logic;
	signal N2_2_39 : std_logic;
	signal N2_3_40 : std_logic;
	signal N2_4_39 : std_logic;
	signal N2_5_40 : std_logic;
	signal N2_6_39 : std_logic;
	signal N2_7_40 : std_logic;
	signal N2_0_40 : std_logic;
	signal N2_1_41 : std_logic;
	signal N2_2_40 : std_logic;
	signal N2_3_41 : std_logic;
	signal N2_4_40 : std_logic;
	signal N2_5_41 : std_logic;
	signal N2_6_40 : std_logic;
	signal N2_7_41 : std_logic;
	signal N2_8_40 : std_logic;
	signal N2_9_41 : std_logic;
	signal N2_0_41 : std_logic;
	signal N2_1_42 : std_logic;
	signal N2_2_41 : std_logic;
	signal N2_3_42 : std_logic;
	signal N2_4_41 : std_logic;
	signal N2_5_42 : std_logic;
	signal N2_6_41 : std_logic;
	signal N2_7_42 : std_logic;
	signal N2_8_41 : std_logic;
	signal N2_9_42 : std_logic;
	signal N2_10_41 : std_logic;
	signal N2_11_42 : std_logic;
	signal N2_0_42 : std_logic;
	signal N2_1_43 : std_logic;
	signal N2_2_42 : std_logic;
	signal N2_3_43 : std_logic;
	signal N2_4_42 : std_logic;
	signal N2_5_43 : std_logic;
	signal N2_6_42 : std_logic;
	signal N2_7_43 : std_logic;
	signal N2_8_42 : std_logic;
	signal N2_9_43 : std_logic;
	signal N2_10_42 : std_logic;
	signal N2_11_43 : std_logic;
	signal N2_12_42 : std_logic;
	signal N2_13_43 : std_logic;
	signal N2_0_43 : std_logic;
	signal N2_1_44 : std_logic;
	signal N2_2_43 : std_logic;
	signal N2_3_44 : std_logic;
	signal N2_4_43 : std_logic;
	signal N2_5_44 : std_logic;
	signal N2_6_43 : std_logic;
	signal N2_7_44 : std_logic;
	signal N2_8_43 : std_logic;
	signal N2_9_44 : std_logic;
	signal N2_10_43 : std_logic;
	signal N2_11_44 : std_logic;
	signal N2_12_43 : std_logic;
	signal N2_13_44 : std_logic;
	signal N2_14_43 : std_logic;
	signal N2_15_44 : std_logic;
	signal N2_0_44 : std_logic;
	signal N2_1_45 : std_logic;
	signal N2_2_44 : std_logic;
	signal N2_3_45 : std_logic;
	signal N2_4_44 : std_logic;
	signal N2_5_45 : std_logic;
	signal N2_6_44 : std_logic;
	signal N2_7_45 : std_logic;
	signal N2_8_44 : std_logic;
	signal N2_9_45 : std_logic;
	signal N2_10_44 : std_logic;
	signal N2_11_45 : std_logic;
	signal N2_12_44 : std_logic;
	signal N2_13_45 : std_logic;
	signal N2_14_44 : std_logic;
	signal N2_15_45 : std_logic;
	signal N2_16_44 : std_logic;
	signal N2_17_45 : std_logic;
	signal N2_0_45 : std_logic;
	signal N2_1_46 : std_logic;
	signal N2_2_45 : std_logic;
	signal N2_3_46 : std_logic;
	signal N2_4_45 : std_logic;
	signal N2_5_46 : std_logic;
	signal N2_6_45 : std_logic;
	signal N2_7_46 : std_logic;
	signal N2_8_45 : std_logic;
	signal N2_9_46 : std_logic;
	signal N2_10_45 : std_logic;
	signal N2_11_46 : std_logic;
	signal N2_12_45 : std_logic;
	signal N2_13_46 : std_logic;
	signal N2_14_45 : std_logic;
	signal N2_15_46 : std_logic;
	signal N2_16_45 : std_logic;
	signal N2_17_46 : std_logic;
	signal N2_18_45 : std_logic;
	signal N2_19_46 : std_logic;
	signal N2_0_46 : std_logic;
	signal N2_1_47 : std_logic;
	signal N2_2_46 : std_logic;
	signal N2_3_47 : std_logic;
	signal N2_4_46 : std_logic;
	signal N2_5_47 : std_logic;
	signal N2_6_46 : std_logic;
	signal N2_7_47 : std_logic;
	signal N2_8_46 : std_logic;
	signal N2_9_47 : std_logic;
	signal N2_10_46 : std_logic;
	signal N2_11_47 : std_logic;
	signal N2_12_46 : std_logic;
	signal N2_13_47 : std_logic;
	signal N2_14_46 : std_logic;
	signal N2_15_47 : std_logic;
	signal N2_16_46 : std_logic;
	signal N2_17_47 : std_logic;
	signal N2_18_46 : std_logic;
	signal N2_19_47 : std_logic;
	signal N2_20_46 : std_logic;
	signal N2_21_47 : std_logic;
	signal N2_0_47 : std_logic;
	signal N2_1_48 : std_logic;
	signal N2_2_47 : std_logic;
	signal N2_3_48 : std_logic;
	signal N2_4_47 : std_logic;
	signal N2_5_48 : std_logic;
	signal N2_6_47 : std_logic;
	signal N2_7_48 : std_logic;
	signal N2_8_47 : std_logic;
	signal N2_9_48 : std_logic;
	signal N2_10_47 : std_logic;
	signal N2_11_48 : std_logic;
	signal N2_12_47 : std_logic;
	signal N2_13_48 : std_logic;
	signal N2_14_47 : std_logic;
	signal N2_15_48 : std_logic;
	signal N2_16_47 : std_logic;
	signal N2_17_48 : std_logic;
	signal N2_18_47 : std_logic;
	signal N2_19_48 : std_logic;
	signal N2_20_47 : std_logic;
	signal N2_21_48 : std_logic;
	signal N2_22_47 : std_logic;
	signal N2_23_48 : std_logic;
	signal N2_0_48 : std_logic;
	signal N2_1_49 : std_logic;
	signal N2_2_48 : std_logic;
	signal N2_3_49 : std_logic;
	signal N2_4_48 : std_logic;
	signal N2_5_49 : std_logic;
	signal N2_6_48 : std_logic;
	signal N2_7_49 : std_logic;
	signal N2_8_48 : std_logic;
	signal N2_9_49 : std_logic;
	signal N2_10_48 : std_logic;
	signal N2_11_49 : std_logic;
	signal N2_12_48 : std_logic;
	signal N2_13_49 : std_logic;
	signal N2_14_48 : std_logic;
	signal N2_15_49 : std_logic;
	signal N2_16_48 : std_logic;
	signal N2_17_49 : std_logic;
	signal N2_18_48 : std_logic;
	signal N2_19_49 : std_logic;
	signal N2_20_48 : std_logic;
	signal N2_21_49 : std_logic;
	signal N2_22_48 : std_logic;
	signal N2_23_49 : std_logic;
	signal N2_24_48 : std_logic;
	signal N2_25_49 : std_logic;
	signal N2_0_49 : std_logic;
	signal N2_1_50 : std_logic;
	signal N2_2_49 : std_logic;
	signal N2_3_50 : std_logic;
	signal N2_4_49 : std_logic;
	signal N2_5_50 : std_logic;
	signal N2_6_49 : std_logic;
	signal N2_7_50 : std_logic;
	signal N2_8_49 : std_logic;
	signal N2_9_50 : std_logic;
	signal N2_10_49 : std_logic;
	signal N2_11_50 : std_logic;
	signal N2_12_49 : std_logic;
	signal N2_13_50 : std_logic;
	signal N2_14_49 : std_logic;
	signal N2_15_50 : std_logic;
	signal N2_16_49 : std_logic;
	signal N2_17_50 : std_logic;
	signal N2_18_49 : std_logic;
	signal N2_19_50 : std_logic;
	signal N2_20_49 : std_logic;
	signal N2_21_50 : std_logic;
	signal N2_22_49 : std_logic;
	signal N2_23_50 : std_logic;
	signal N2_24_49 : std_logic;
	signal N2_25_50 : std_logic;
	signal N2_26_49 : std_logic;
	signal N2_27_50 : std_logic;
	signal N2_0_50 : std_logic;
	signal N2_1_51 : std_logic;
	signal N2_2_50 : std_logic;
	signal N2_3_51 : std_logic;
	signal N2_4_50 : std_logic;
	signal N2_5_51 : std_logic;
	signal N2_6_50 : std_logic;
	signal N2_7_51 : std_logic;
	signal N2_8_50 : std_logic;
	signal N2_9_51 : std_logic;
	signal N2_10_50 : std_logic;
	signal N2_11_51 : std_logic;
	signal N2_12_50 : std_logic;
	signal N2_13_51 : std_logic;
	signal N2_14_50 : std_logic;
	signal N2_15_51 : std_logic;
	signal N2_16_50 : std_logic;
	signal N2_17_51 : std_logic;
	signal N2_18_50 : std_logic;
	signal N2_19_51 : std_logic;
	signal N2_20_50 : std_logic;
	signal N2_21_51 : std_logic;
	signal N2_22_50 : std_logic;
	signal N2_23_51 : std_logic;
	signal N2_24_50 : std_logic;
	signal N2_25_51 : std_logic;
	signal N2_26_50 : std_logic;
	signal N2_27_51 : std_logic;
	signal N2_28_50 : std_logic;
	signal N2_29_51 : std_logic;
	signal N2_0_51 : std_logic;
	signal N2_1_52 : std_logic;
	signal N2_2_51 : std_logic;
	signal N2_3_52 : std_logic;
	signal N2_4_51 : std_logic;
	signal N2_5_52 : std_logic;
	signal N2_6_51 : std_logic;
	signal N2_7_52 : std_logic;
	signal N2_8_51 : std_logic;
	signal N2_9_52 : std_logic;
	signal N2_10_51 : std_logic;
	signal N2_11_52 : std_logic;
	signal N2_12_51 : std_logic;
	signal N2_13_52 : std_logic;
	signal N2_14_51 : std_logic;
	signal N2_15_52 : std_logic;
	signal N2_16_51 : std_logic;
	signal N2_17_52 : std_logic;
	signal N2_18_51 : std_logic;
	signal N2_19_52 : std_logic;
	signal N2_20_51 : std_logic;
	signal N2_21_52 : std_logic;
	signal N2_22_51 : std_logic;
	signal N2_23_52 : std_logic;
	signal N2_24_51 : std_logic;
	signal N2_25_52 : std_logic;
	signal N2_26_51 : std_logic;
	signal N2_27_52 : std_logic;
	signal N2_28_51 : std_logic;
	signal N2_29_52 : std_logic;
	signal N2_30_51 : std_logic;
	signal N2_31_52 : std_logic;
	signal N2_0_52 : std_logic;
	signal N2_1_53 : std_logic;
	signal N2_2_52 : std_logic;
	signal N2_3_53 : std_logic;
	signal N2_4_52 : std_logic;
	signal N2_5_53 : std_logic;
	signal N2_6_52 : std_logic;
	signal N2_7_53 : std_logic;
	signal N2_8_52 : std_logic;
	signal N2_9_53 : std_logic;
	signal N2_10_52 : std_logic;
	signal N2_11_53 : std_logic;
	signal N2_12_52 : std_logic;
	signal N2_13_53 : std_logic;
	signal N2_14_52 : std_logic;
	signal N2_15_53 : std_logic;
	signal N2_16_52 : std_logic;
	signal N2_17_53 : std_logic;
	signal N2_18_52 : std_logic;
	signal N2_19_53 : std_logic;
	signal N2_20_52 : std_logic;
	signal N2_21_53 : std_logic;
	signal N2_22_52 : std_logic;
	signal N2_23_53 : std_logic;
	signal N2_24_52 : std_logic;
	signal N2_25_53 : std_logic;
	signal N2_26_52 : std_logic;
	signal N2_27_53 : std_logic;
	signal N2_28_52 : std_logic;
	signal N2_29_53 : std_logic;
	signal N2_30_52 : std_logic;
	signal N2_31_53 : std_logic;
	signal N2_32_52 : std_logic;
	signal N2_33_53 : std_logic;
	signal N2_0_53 : std_logic;
	signal N2_1_54 : std_logic;
	signal N2_2_53 : std_logic;
	signal N2_3_54 : std_logic;
	signal N2_4_53 : std_logic;
	signal N2_5_54 : std_logic;
	signal N2_6_53 : std_logic;
	signal N2_7_54 : std_logic;
	signal N2_8_53 : std_logic;
	signal N2_9_54 : std_logic;
	signal N2_10_53 : std_logic;
	signal N2_11_54 : std_logic;
	signal N2_12_53 : std_logic;
	signal N2_13_54 : std_logic;
	signal N2_14_53 : std_logic;
	signal N2_15_54 : std_logic;
	signal N2_16_53 : std_logic;
	signal N2_17_54 : std_logic;
	signal N2_18_53 : std_logic;
	signal N2_19_54 : std_logic;
	signal N2_20_53 : std_logic;
	signal N2_21_54 : std_logic;
	signal N2_22_53 : std_logic;
	signal N2_23_54 : std_logic;
	signal N2_24_53 : std_logic;
	signal N2_25_54 : std_logic;
	signal N2_26_53 : std_logic;
	signal N2_27_54 : std_logic;
	signal N2_28_53 : std_logic;
	signal N2_29_54 : std_logic;
	signal N2_30_53 : std_logic;
	signal N2_31_54 : std_logic;
	signal N2_32_53 : std_logic;
	signal N2_33_54 : std_logic;
	signal N2_0_54 : std_logic;
	signal N2_1_55 : std_logic;
	signal N2_2_54 : std_logic;
	signal N2_3_55 : std_logic;
	signal N2_4_54 : std_logic;
	signal N2_5_55 : std_logic;
	signal N2_6_54 : std_logic;
	signal N2_7_55 : std_logic;
	signal N2_8_54 : std_logic;
	signal N2_9_55 : std_logic;
	signal N2_10_54 : std_logic;
	signal N2_11_55 : std_logic;
	signal N2_12_54 : std_logic;
	signal N2_13_55 : std_logic;
	signal N2_14_54 : std_logic;
	signal N2_15_55 : std_logic;
	signal N2_16_54 : std_logic;
	signal N2_17_55 : std_logic;
	signal N2_18_54 : std_logic;
	signal N2_19_55 : std_logic;
	signal N2_20_54 : std_logic;
	signal N2_21_55 : std_logic;
	signal N2_22_54 : std_logic;
	signal N2_23_55 : std_logic;
	signal N2_24_54 : std_logic;
	signal N2_25_55 : std_logic;
	signal N2_26_54 : std_logic;
	signal N2_27_55 : std_logic;
	signal N2_28_54 : std_logic;
	signal N2_29_55 : std_logic;
	signal N2_30_54 : std_logic;
	signal N2_31_55 : std_logic;
	signal N2_0_55 : std_logic;
	signal N2_1_56 : std_logic;
	signal N2_2_55 : std_logic;
	signal N2_3_56 : std_logic;
	signal N2_4_55 : std_logic;
	signal N2_5_56 : std_logic;
	signal N2_6_55 : std_logic;
	signal N2_7_56 : std_logic;
	signal N2_8_55 : std_logic;
	signal N2_9_56 : std_logic;
	signal N2_10_55 : std_logic;
	signal N2_11_56 : std_logic;
	signal N2_12_55 : std_logic;
	signal N2_13_56 : std_logic;
	signal N2_14_55 : std_logic;
	signal N2_15_56 : std_logic;
	signal N2_16_55 : std_logic;
	signal N2_17_56 : std_logic;
	signal N2_18_55 : std_logic;
	signal N2_19_56 : std_logic;
	signal N2_20_55 : std_logic;
	signal N2_21_56 : std_logic;
	signal N2_22_55 : std_logic;
	signal N2_23_56 : std_logic;
	signal N2_24_55 : std_logic;
	signal N2_25_56 : std_logic;
	signal N2_26_55 : std_logic;
	signal N2_27_56 : std_logic;
	signal N2_28_55 : std_logic;
	signal N2_29_56 : std_logic;
	signal N2_0_56 : std_logic;
	signal N2_1_57 : std_logic;
	signal N2_2_56 : std_logic;
	signal N2_3_57 : std_logic;
	signal N2_4_56 : std_logic;
	signal N2_5_57 : std_logic;
	signal N2_6_56 : std_logic;
	signal N2_7_57 : std_logic;
	signal N2_8_56 : std_logic;
	signal N2_9_57 : std_logic;
	signal N2_10_56 : std_logic;
	signal N2_11_57 : std_logic;
	signal N2_12_56 : std_logic;
	signal N2_13_57 : std_logic;
	signal N2_14_56 : std_logic;
	signal N2_15_57 : std_logic;
	signal N2_16_56 : std_logic;
	signal N2_17_57 : std_logic;
	signal N2_18_56 : std_logic;
	signal N2_19_57 : std_logic;
	signal N2_20_56 : std_logic;
	signal N2_21_57 : std_logic;
	signal N2_22_56 : std_logic;
	signal N2_23_57 : std_logic;
	signal N2_24_56 : std_logic;
	signal N2_25_57 : std_logic;
	signal N2_26_56 : std_logic;
	signal N2_27_57 : std_logic;
	signal N2_0_57 : std_logic;
	signal N2_1_58 : std_logic;
	signal N2_2_57 : std_logic;
	signal N2_3_58 : std_logic;
	signal N2_4_57 : std_logic;
	signal N2_5_58 : std_logic;
	signal N2_6_57 : std_logic;
	signal N2_7_58 : std_logic;
	signal N2_8_57 : std_logic;
	signal N2_9_58 : std_logic;
	signal N2_10_57 : std_logic;
	signal N2_11_58 : std_logic;
	signal N2_12_57 : std_logic;
	signal N2_13_58 : std_logic;
	signal N2_14_57 : std_logic;
	signal N2_15_58 : std_logic;
	signal N2_16_57 : std_logic;
	signal N2_17_58 : std_logic;
	signal N2_18_57 : std_logic;
	signal N2_19_58 : std_logic;
	signal N2_20_57 : std_logic;
	signal N2_21_58 : std_logic;
	signal N2_22_57 : std_logic;
	signal N2_23_58 : std_logic;
	signal N2_24_57 : std_logic;
	signal N2_25_58 : std_logic;
	signal N2_0_58 : std_logic;
	signal N2_1_59 : std_logic;
	signal N2_2_58 : std_logic;
	signal N2_3_59 : std_logic;
	signal N2_4_58 : std_logic;
	signal N2_5_59 : std_logic;
	signal N2_6_58 : std_logic;
	signal N2_7_59 : std_logic;
	signal N2_8_58 : std_logic;
	signal N2_9_59 : std_logic;
	signal N2_10_58 : std_logic;
	signal N2_11_59 : std_logic;
	signal N2_12_58 : std_logic;
	signal N2_13_59 : std_logic;
	signal N2_14_58 : std_logic;
	signal N2_15_59 : std_logic;
	signal N2_16_58 : std_logic;
	signal N2_17_59 : std_logic;
	signal N2_18_58 : std_logic;
	signal N2_19_59 : std_logic;
	signal N2_20_58 : std_logic;
	signal N2_21_59 : std_logic;
	signal N2_22_58 : std_logic;
	signal N2_23_59 : std_logic;
	signal N2_0_59 : std_logic;
	signal N2_1_60 : std_logic;
	signal N2_2_59 : std_logic;
	signal N2_3_60 : std_logic;
	signal N2_4_59 : std_logic;
	signal N2_5_60 : std_logic;
	signal N2_6_59 : std_logic;
	signal N2_7_60 : std_logic;
	signal N2_8_59 : std_logic;
	signal N2_9_60 : std_logic;
	signal N2_10_59 : std_logic;
	signal N2_11_60 : std_logic;
	signal N2_12_59 : std_logic;
	signal N2_13_60 : std_logic;
	signal N2_14_59 : std_logic;
	signal N2_15_60 : std_logic;
	signal N2_16_59 : std_logic;
	signal N2_17_60 : std_logic;
	signal N2_18_59 : std_logic;
	signal N2_19_60 : std_logic;
	signal N2_20_59 : std_logic;
	signal N2_21_60 : std_logic;
	signal N2_0_60 : std_logic;
	signal N2_1_61 : std_logic;
	signal N2_2_60 : std_logic;
	signal N2_3_61 : std_logic;
	signal N2_4_60 : std_logic;
	signal N2_5_61 : std_logic;
	signal N2_6_60 : std_logic;
	signal N2_7_61 : std_logic;
	signal N2_8_60 : std_logic;
	signal N2_9_61 : std_logic;
	signal N2_10_60 : std_logic;
	signal N2_11_61 : std_logic;
	signal N2_12_60 : std_logic;
	signal N2_13_61 : std_logic;
	signal N2_14_60 : std_logic;
	signal N2_15_61 : std_logic;
	signal N2_16_60 : std_logic;
	signal N2_17_61 : std_logic;
	signal N2_18_60 : std_logic;
	signal N2_19_61 : std_logic;
	signal N2_0_61 : std_logic;
	signal N2_1_62 : std_logic;
	signal N2_2_61 : std_logic;
	signal N2_3_62 : std_logic;
	signal N2_4_61 : std_logic;
	signal N2_5_62 : std_logic;
	signal N2_6_61 : std_logic;
	signal N2_7_62 : std_logic;
	signal N2_8_61 : std_logic;
	signal N2_9_62 : std_logic;
	signal N2_10_61 : std_logic;
	signal N2_11_62 : std_logic;
	signal N2_12_61 : std_logic;
	signal N2_13_62 : std_logic;
	signal N2_14_61 : std_logic;
	signal N2_15_62 : std_logic;
	signal N2_16_61 : std_logic;
	signal N2_17_62 : std_logic;
	signal N2_0_62 : std_logic;
	signal N2_1_63 : std_logic;
	signal N2_2_62 : std_logic;
	signal N2_3_63 : std_logic;
	signal N2_4_62 : std_logic;
	signal N2_5_63 : std_logic;
	signal N2_6_62 : std_logic;
	signal N2_7_63 : std_logic;
	signal N2_8_62 : std_logic;
	signal N2_9_63 : std_logic;
	signal N2_10_62 : std_logic;
	signal N2_11_63 : std_logic;
	signal N2_12_62 : std_logic;
	signal N2_13_63 : std_logic;
	signal N2_14_62 : std_logic;
	signal N2_15_63 : std_logic;
	signal N2_0_63 : std_logic;
	signal N2_1_64 : std_logic;
	signal N2_2_63 : std_logic;
	signal N2_3_64 : std_logic;
	signal N2_4_63 : std_logic;
	signal N2_5_64 : std_logic;
	signal N2_6_63 : std_logic;
	signal N2_7_64 : std_logic;
	signal N2_8_63 : std_logic;
	signal N2_9_64 : std_logic;
	signal N2_10_63 : std_logic;
	signal N2_11_64 : std_logic;
	signal N2_12_63 : std_logic;
	signal N2_13_64 : std_logic;
	signal N2_0_64 : std_logic;
	signal N2_1_65 : std_logic;
	signal N2_2_64 : std_logic;
	signal N2_3_65 : std_logic;
	signal N2_4_64 : std_logic;
	signal N2_5_65 : std_logic;
	signal N2_6_64 : std_logic;
	signal N2_7_65 : std_logic;
	signal N2_8_64 : std_logic;
	signal N2_9_65 : std_logic;
	signal N2_10_64 : std_logic;
	signal N2_11_65 : std_logic;
	signal N2_0_65 : std_logic;
	signal N2_1_66 : std_logic;
	signal N2_2_65 : std_logic;
	signal N2_3_66 : std_logic;
	signal N2_4_65 : std_logic;
	signal N2_5_66 : std_logic;
	signal N2_6_65 : std_logic;
	signal N2_7_66 : std_logic;
	signal N2_8_65 : std_logic;
	signal N2_9_66 : std_logic;
	signal N2_0_66 : std_logic;
	signal N2_1_67 : std_logic;
	signal N2_2_66 : std_logic;
	signal N2_3_67 : std_logic;
	signal N2_4_66 : std_logic;
	signal N2_5_67 : std_logic;
	signal N2_6_66 : std_logic;
	signal N2_7_67 : std_logic;
	signal N2_0_67 : std_logic;
	signal N2_1_68 : std_logic;
	signal N2_2_67 : std_logic;
	signal N2_3_68 : std_logic;
	signal N2_4_67 : std_logic;
	signal N2_5_68 : std_logic;
	signal N2_0_68 : std_logic;
	signal N2_1_69 : std_logic;
	signal N2_2_68 : std_logic;
	signal N2_3_69 : std_logic;
	signal N2_0_69 : std_logic;
	signal N2_1_70 : std_logic;
	signal N3_0_24 : std_logic;
	signal N3_1_25 : std_logic;
	signal N3_0_25 : std_logic;
	signal N3_1_26 : std_logic;
	signal N3_2_25 : std_logic;
	signal N3_3_26 : std_logic;
	signal N3_0_26 : std_logic;
	signal N3_1_27 : std_logic;
	signal N3_2_26 : std_logic;
	signal N3_3_27 : std_logic;
	signal N3_4_26 : std_logic;
	signal N3_5_27 : std_logic;
	signal N3_0_27 : std_logic;
	signal N3_1_28 : std_logic;
	signal N3_2_27 : std_logic;
	signal N3_3_28 : std_logic;
	signal N3_4_27 : std_logic;
	signal N3_5_28 : std_logic;
	signal N3_6_27 : std_logic;
	signal N3_7_28 : std_logic;
	signal N3_0_28 : std_logic;
	signal N3_1_29 : std_logic;
	signal N3_2_28 : std_logic;
	signal N3_3_29 : std_logic;
	signal N3_4_28 : std_logic;
	signal N3_5_29 : std_logic;
	signal N3_6_28 : std_logic;
	signal N3_7_29 : std_logic;
	signal N3_8_28 : std_logic;
	signal N3_9_29 : std_logic;
	signal N3_0_29 : std_logic;
	signal N3_1_30 : std_logic;
	signal N3_2_29 : std_logic;
	signal N3_3_30 : std_logic;
	signal N3_4_29 : std_logic;
	signal N3_5_30 : std_logic;
	signal N3_6_29 : std_logic;
	signal N3_7_30 : std_logic;
	signal N3_8_29 : std_logic;
	signal N3_9_30 : std_logic;
	signal N3_10_29 : std_logic;
	signal N3_11_30 : std_logic;
	signal N3_0_30 : std_logic;
	signal N3_1_31 : std_logic;
	signal N3_2_30 : std_logic;
	signal N3_3_31 : std_logic;
	signal N3_4_30 : std_logic;
	signal N3_5_31 : std_logic;
	signal N3_6_30 : std_logic;
	signal N3_7_31 : std_logic;
	signal N3_8_30 : std_logic;
	signal N3_9_31 : std_logic;
	signal N3_10_30 : std_logic;
	signal N3_11_31 : std_logic;
	signal N3_12_30 : std_logic;
	signal N3_13_31 : std_logic;
	signal N3_0_31 : std_logic;
	signal N3_1_32 : std_logic;
	signal N3_2_31 : std_logic;
	signal N3_3_32 : std_logic;
	signal N3_4_31 : std_logic;
	signal N3_5_32 : std_logic;
	signal N3_6_31 : std_logic;
	signal N3_7_32 : std_logic;
	signal N3_8_31 : std_logic;
	signal N3_9_32 : std_logic;
	signal N3_10_31 : std_logic;
	signal N3_11_32 : std_logic;
	signal N3_12_31 : std_logic;
	signal N3_13_32 : std_logic;
	signal N3_14_31 : std_logic;
	signal N3_15_32 : std_logic;
	signal N3_0_32 : std_logic;
	signal N3_1_33 : std_logic;
	signal N3_2_32 : std_logic;
	signal N3_3_33 : std_logic;
	signal N3_4_32 : std_logic;
	signal N3_5_33 : std_logic;
	signal N3_6_32 : std_logic;
	signal N3_7_33 : std_logic;
	signal N3_8_32 : std_logic;
	signal N3_9_33 : std_logic;
	signal N3_10_32 : std_logic;
	signal N3_11_33 : std_logic;
	signal N3_12_32 : std_logic;
	signal N3_13_33 : std_logic;
	signal N3_14_32 : std_logic;
	signal N3_15_33 : std_logic;
	signal N3_16_32 : std_logic;
	signal N3_17_33 : std_logic;
	signal N3_0_33 : std_logic;
	signal N3_1_34 : std_logic;
	signal N3_2_33 : std_logic;
	signal N3_3_34 : std_logic;
	signal N3_4_33 : std_logic;
	signal N3_5_34 : std_logic;
	signal N3_6_33 : std_logic;
	signal N3_7_34 : std_logic;
	signal N3_8_33 : std_logic;
	signal N3_9_34 : std_logic;
	signal N3_10_33 : std_logic;
	signal N3_11_34 : std_logic;
	signal N3_12_33 : std_logic;
	signal N3_13_34 : std_logic;
	signal N3_14_33 : std_logic;
	signal N3_15_34 : std_logic;
	signal N3_16_33 : std_logic;
	signal N3_17_34 : std_logic;
	signal N3_18_33 : std_logic;
	signal N3_19_34 : std_logic;
	signal N3_0_34 : std_logic;
	signal N3_1_35 : std_logic;
	signal N3_2_34 : std_logic;
	signal N3_3_35 : std_logic;
	signal N3_4_34 : std_logic;
	signal N3_5_35 : std_logic;
	signal N3_6_34 : std_logic;
	signal N3_7_35 : std_logic;
	signal N3_8_34 : std_logic;
	signal N3_9_35 : std_logic;
	signal N3_10_34 : std_logic;
	signal N3_11_35 : std_logic;
	signal N3_12_34 : std_logic;
	signal N3_13_35 : std_logic;
	signal N3_14_34 : std_logic;
	signal N3_15_35 : std_logic;
	signal N3_16_34 : std_logic;
	signal N3_17_35 : std_logic;
	signal N3_18_34 : std_logic;
	signal N3_19_35 : std_logic;
	signal N3_20_34 : std_logic;
	signal N3_21_35 : std_logic;
	signal N3_0_35 : std_logic;
	signal N3_1_36 : std_logic;
	signal N3_2_35 : std_logic;
	signal N3_3_36 : std_logic;
	signal N3_4_35 : std_logic;
	signal N3_5_36 : std_logic;
	signal N3_6_35 : std_logic;
	signal N3_7_36 : std_logic;
	signal N3_8_35 : std_logic;
	signal N3_9_36 : std_logic;
	signal N3_10_35 : std_logic;
	signal N3_11_36 : std_logic;
	signal N3_12_35 : std_logic;
	signal N3_13_36 : std_logic;
	signal N3_14_35 : std_logic;
	signal N3_15_36 : std_logic;
	signal N3_16_35 : std_logic;
	signal N3_17_36 : std_logic;
	signal N3_18_35 : std_logic;
	signal N3_19_36 : std_logic;
	signal N3_20_35 : std_logic;
	signal N3_21_36 : std_logic;
	signal N3_22_35 : std_logic;
	signal N3_23_36 : std_logic;
	signal N3_0_36 : std_logic;
	signal N3_1_37 : std_logic;
	signal N3_2_36 : std_logic;
	signal N3_3_37 : std_logic;
	signal N3_4_36 : std_logic;
	signal N3_5_37 : std_logic;
	signal N3_6_36 : std_logic;
	signal N3_7_37 : std_logic;
	signal N3_8_36 : std_logic;
	signal N3_9_37 : std_logic;
	signal N3_10_36 : std_logic;
	signal N3_11_37 : std_logic;
	signal N3_12_36 : std_logic;
	signal N3_13_37 : std_logic;
	signal N3_14_36 : std_logic;
	signal N3_15_37 : std_logic;
	signal N3_16_36 : std_logic;
	signal N3_17_37 : std_logic;
	signal N3_18_36 : std_logic;
	signal N3_19_37 : std_logic;
	signal N3_20_36 : std_logic;
	signal N3_21_37 : std_logic;
	signal N3_22_36 : std_logic;
	signal N3_23_37 : std_logic;
	signal N3_0_37 : std_logic;
	signal N3_1_38 : std_logic;
	signal N3_2_37 : std_logic;
	signal N3_3_38 : std_logic;
	signal N3_4_37 : std_logic;
	signal N3_5_38 : std_logic;
	signal N3_6_37 : std_logic;
	signal N3_7_38 : std_logic;
	signal N3_8_37 : std_logic;
	signal N3_9_38 : std_logic;
	signal N3_10_37 : std_logic;
	signal N3_11_38 : std_logic;
	signal N3_12_37 : std_logic;
	signal N3_13_38 : std_logic;
	signal N3_14_37 : std_logic;
	signal N3_15_38 : std_logic;
	signal N3_16_37 : std_logic;
	signal N3_17_38 : std_logic;
	signal N3_18_37 : std_logic;
	signal N3_19_38 : std_logic;
	signal N3_20_37 : std_logic;
	signal N3_21_38 : std_logic;
	signal N3_22_37 : std_logic;
	signal N3_23_38 : std_logic;
	signal N3_0_38 : std_logic;
	signal N3_1_39 : std_logic;
	signal N3_2_38 : std_logic;
	signal N3_3_39 : std_logic;
	signal N3_4_38 : std_logic;
	signal N3_5_39 : std_logic;
	signal N3_6_38 : std_logic;
	signal N3_7_39 : std_logic;
	signal N3_8_38 : std_logic;
	signal N3_9_39 : std_logic;
	signal N3_10_38 : std_logic;
	signal N3_11_39 : std_logic;
	signal N3_12_38 : std_logic;
	signal N3_13_39 : std_logic;
	signal N3_14_38 : std_logic;
	signal N3_15_39 : std_logic;
	signal N3_16_38 : std_logic;
	signal N3_17_39 : std_logic;
	signal N3_18_38 : std_logic;
	signal N3_19_39 : std_logic;
	signal N3_20_38 : std_logic;
	signal N3_21_39 : std_logic;
	signal N3_22_38 : std_logic;
	signal N3_23_39 : std_logic;
	signal N3_0_39 : std_logic;
	signal N3_1_40 : std_logic;
	signal N3_2_39 : std_logic;
	signal N3_3_40 : std_logic;
	signal N3_4_39 : std_logic;
	signal N3_5_40 : std_logic;
	signal N3_6_39 : std_logic;
	signal N3_7_40 : std_logic;
	signal N3_8_39 : std_logic;
	signal N3_9_40 : std_logic;
	signal N3_10_39 : std_logic;
	signal N3_11_40 : std_logic;
	signal N3_12_39 : std_logic;
	signal N3_13_40 : std_logic;
	signal N3_14_39 : std_logic;
	signal N3_15_40 : std_logic;
	signal N3_16_39 : std_logic;
	signal N3_17_40 : std_logic;
	signal N3_18_39 : std_logic;
	signal N3_19_40 : std_logic;
	signal N3_20_39 : std_logic;
	signal N3_21_40 : std_logic;
	signal N3_22_39 : std_logic;
	signal N3_23_40 : std_logic;
	signal N3_0_40 : std_logic;
	signal N3_1_41 : std_logic;
	signal N3_2_40 : std_logic;
	signal N3_3_41 : std_logic;
	signal N3_4_40 : std_logic;
	signal N3_5_41 : std_logic;
	signal N3_6_40 : std_logic;
	signal N3_7_41 : std_logic;
	signal N3_8_40 : std_logic;
	signal N3_9_41 : std_logic;
	signal N3_10_40 : std_logic;
	signal N3_11_41 : std_logic;
	signal N3_12_40 : std_logic;
	signal N3_13_41 : std_logic;
	signal N3_14_40 : std_logic;
	signal N3_15_41 : std_logic;
	signal N3_16_40 : std_logic;
	signal N3_17_41 : std_logic;
	signal N3_18_40 : std_logic;
	signal N3_19_41 : std_logic;
	signal N3_20_40 : std_logic;
	signal N3_21_41 : std_logic;
	signal N3_22_40 : std_logic;
	signal N3_23_41 : std_logic;
	signal N3_0_41 : std_logic;
	signal N3_1_42 : std_logic;
	signal N3_2_41 : std_logic;
	signal N3_3_42 : std_logic;
	signal N3_4_41 : std_logic;
	signal N3_5_42 : std_logic;
	signal N3_6_41 : std_logic;
	signal N3_7_42 : std_logic;
	signal N3_8_41 : std_logic;
	signal N3_9_42 : std_logic;
	signal N3_10_41 : std_logic;
	signal N3_11_42 : std_logic;
	signal N3_12_41 : std_logic;
	signal N3_13_42 : std_logic;
	signal N3_14_41 : std_logic;
	signal N3_15_42 : std_logic;
	signal N3_16_41 : std_logic;
	signal N3_17_42 : std_logic;
	signal N3_18_41 : std_logic;
	signal N3_19_42 : std_logic;
	signal N3_20_41 : std_logic;
	signal N3_21_42 : std_logic;
	signal N3_22_41 : std_logic;
	signal N3_23_42 : std_logic;
	signal N3_0_42 : std_logic;
	signal N3_1_43 : std_logic;
	signal N3_2_42 : std_logic;
	signal N3_3_43 : std_logic;
	signal N3_4_42 : std_logic;
	signal N3_5_43 : std_logic;
	signal N3_6_42 : std_logic;
	signal N3_7_43 : std_logic;
	signal N3_8_42 : std_logic;
	signal N3_9_43 : std_logic;
	signal N3_10_42 : std_logic;
	signal N3_11_43 : std_logic;
	signal N3_12_42 : std_logic;
	signal N3_13_43 : std_logic;
	signal N3_14_42 : std_logic;
	signal N3_15_43 : std_logic;
	signal N3_16_42 : std_logic;
	signal N3_17_43 : std_logic;
	signal N3_18_42 : std_logic;
	signal N3_19_43 : std_logic;
	signal N3_20_42 : std_logic;
	signal N3_21_43 : std_logic;
	signal N3_22_42 : std_logic;
	signal N3_23_43 : std_logic;
	signal N3_0_43 : std_logic;
	signal N3_1_44 : std_logic;
	signal N3_2_43 : std_logic;
	signal N3_3_44 : std_logic;
	signal N3_4_43 : std_logic;
	signal N3_5_44 : std_logic;
	signal N3_6_43 : std_logic;
	signal N3_7_44 : std_logic;
	signal N3_8_43 : std_logic;
	signal N3_9_44 : std_logic;
	signal N3_10_43 : std_logic;
	signal N3_11_44 : std_logic;
	signal N3_12_43 : std_logic;
	signal N3_13_44 : std_logic;
	signal N3_14_43 : std_logic;
	signal N3_15_44 : std_logic;
	signal N3_16_43 : std_logic;
	signal N3_17_44 : std_logic;
	signal N3_18_43 : std_logic;
	signal N3_19_44 : std_logic;
	signal N3_20_43 : std_logic;
	signal N3_21_44 : std_logic;
	signal N3_22_43 : std_logic;
	signal N3_23_44 : std_logic;
	signal N3_0_44 : std_logic;
	signal N3_1_45 : std_logic;
	signal N3_2_44 : std_logic;
	signal N3_3_45 : std_logic;
	signal N3_4_44 : std_logic;
	signal N3_5_45 : std_logic;
	signal N3_6_44 : std_logic;
	signal N3_7_45 : std_logic;
	signal N3_8_44 : std_logic;
	signal N3_9_45 : std_logic;
	signal N3_10_44 : std_logic;
	signal N3_11_45 : std_logic;
	signal N3_12_44 : std_logic;
	signal N3_13_45 : std_logic;
	signal N3_14_44 : std_logic;
	signal N3_15_45 : std_logic;
	signal N3_16_44 : std_logic;
	signal N3_17_45 : std_logic;
	signal N3_18_44 : std_logic;
	signal N3_19_45 : std_logic;
	signal N3_20_44 : std_logic;
	signal N3_21_45 : std_logic;
	signal N3_22_44 : std_logic;
	signal N3_23_45 : std_logic;
	signal N3_0_45 : std_logic;
	signal N3_1_46 : std_logic;
	signal N3_2_45 : std_logic;
	signal N3_3_46 : std_logic;
	signal N3_4_45 : std_logic;
	signal N3_5_46 : std_logic;
	signal N3_6_45 : std_logic;
	signal N3_7_46 : std_logic;
	signal N3_8_45 : std_logic;
	signal N3_9_46 : std_logic;
	signal N3_10_45 : std_logic;
	signal N3_11_46 : std_logic;
	signal N3_12_45 : std_logic;
	signal N3_13_46 : std_logic;
	signal N3_14_45 : std_logic;
	signal N3_15_46 : std_logic;
	signal N3_16_45 : std_logic;
	signal N3_17_46 : std_logic;
	signal N3_18_45 : std_logic;
	signal N3_19_46 : std_logic;
	signal N3_20_45 : std_logic;
	signal N3_21_46 : std_logic;
	signal N3_22_45 : std_logic;
	signal N3_23_46 : std_logic;
	signal N3_0_46 : std_logic;
	signal N3_1_47 : std_logic;
	signal N3_2_46 : std_logic;
	signal N3_3_47 : std_logic;
	signal N3_4_46 : std_logic;
	signal N3_5_47 : std_logic;
	signal N3_6_46 : std_logic;
	signal N3_7_47 : std_logic;
	signal N3_8_46 : std_logic;
	signal N3_9_47 : std_logic;
	signal N3_10_46 : std_logic;
	signal N3_11_47 : std_logic;
	signal N3_12_46 : std_logic;
	signal N3_13_47 : std_logic;
	signal N3_14_46 : std_logic;
	signal N3_15_47 : std_logic;
	signal N3_16_46 : std_logic;
	signal N3_17_47 : std_logic;
	signal N3_18_46 : std_logic;
	signal N3_19_47 : std_logic;
	signal N3_20_46 : std_logic;
	signal N3_21_47 : std_logic;
	signal N3_22_46 : std_logic;
	signal N3_23_47 : std_logic;
	signal N3_0_47 : std_logic;
	signal N3_1_48 : std_logic;
	signal N3_2_47 : std_logic;
	signal N3_3_48 : std_logic;
	signal N3_4_47 : std_logic;
	signal N3_5_48 : std_logic;
	signal N3_6_47 : std_logic;
	signal N3_7_48 : std_logic;
	signal N3_8_47 : std_logic;
	signal N3_9_48 : std_logic;
	signal N3_10_47 : std_logic;
	signal N3_11_48 : std_logic;
	signal N3_12_47 : std_logic;
	signal N3_13_48 : std_logic;
	signal N3_14_47 : std_logic;
	signal N3_15_48 : std_logic;
	signal N3_16_47 : std_logic;
	signal N3_17_48 : std_logic;
	signal N3_18_47 : std_logic;
	signal N3_19_48 : std_logic;
	signal N3_20_47 : std_logic;
	signal N3_21_48 : std_logic;
	signal N3_22_47 : std_logic;
	signal N3_23_48 : std_logic;
	signal N3_0_48 : std_logic;
	signal N3_1_49 : std_logic;
	signal N3_2_48 : std_logic;
	signal N3_3_49 : std_logic;
	signal N3_4_48 : std_logic;
	signal N3_5_49 : std_logic;
	signal N3_6_48 : std_logic;
	signal N3_7_49 : std_logic;
	signal N3_8_48 : std_logic;
	signal N3_9_49 : std_logic;
	signal N3_10_48 : std_logic;
	signal N3_11_49 : std_logic;
	signal N3_12_48 : std_logic;
	signal N3_13_49 : std_logic;
	signal N3_14_48 : std_logic;
	signal N3_15_49 : std_logic;
	signal N3_16_48 : std_logic;
	signal N3_17_49 : std_logic;
	signal N3_18_48 : std_logic;
	signal N3_19_49 : std_logic;
	signal N3_20_48 : std_logic;
	signal N3_21_49 : std_logic;
	signal N3_22_48 : std_logic;
	signal N3_23_49 : std_logic;
	signal N3_0_49 : std_logic;
	signal N3_1_50 : std_logic;
	signal N3_2_49 : std_logic;
	signal N3_3_50 : std_logic;
	signal N3_4_49 : std_logic;
	signal N3_5_50 : std_logic;
	signal N3_6_49 : std_logic;
	signal N3_7_50 : std_logic;
	signal N3_8_49 : std_logic;
	signal N3_9_50 : std_logic;
	signal N3_10_49 : std_logic;
	signal N3_11_50 : std_logic;
	signal N3_12_49 : std_logic;
	signal N3_13_50 : std_logic;
	signal N3_14_49 : std_logic;
	signal N3_15_50 : std_logic;
	signal N3_16_49 : std_logic;
	signal N3_17_50 : std_logic;
	signal N3_18_49 : std_logic;
	signal N3_19_50 : std_logic;
	signal N3_20_49 : std_logic;
	signal N3_21_50 : std_logic;
	signal N3_22_49 : std_logic;
	signal N3_23_50 : std_logic;
	signal N3_0_50 : std_logic;
	signal N3_1_51 : std_logic;
	signal N3_2_50 : std_logic;
	signal N3_3_51 : std_logic;
	signal N3_4_50 : std_logic;
	signal N3_5_51 : std_logic;
	signal N3_6_50 : std_logic;
	signal N3_7_51 : std_logic;
	signal N3_8_50 : std_logic;
	signal N3_9_51 : std_logic;
	signal N3_10_50 : std_logic;
	signal N3_11_51 : std_logic;
	signal N3_12_50 : std_logic;
	signal N3_13_51 : std_logic;
	signal N3_14_50 : std_logic;
	signal N3_15_51 : std_logic;
	signal N3_16_50 : std_logic;
	signal N3_17_51 : std_logic;
	signal N3_18_50 : std_logic;
	signal N3_19_51 : std_logic;
	signal N3_20_50 : std_logic;
	signal N3_21_51 : std_logic;
	signal N3_22_50 : std_logic;
	signal N3_23_51 : std_logic;
	signal N3_0_51 : std_logic;
	signal N3_1_52 : std_logic;
	signal N3_2_51 : std_logic;
	signal N3_3_52 : std_logic;
	signal N3_4_51 : std_logic;
	signal N3_5_52 : std_logic;
	signal N3_6_51 : std_logic;
	signal N3_7_52 : std_logic;
	signal N3_8_51 : std_logic;
	signal N3_9_52 : std_logic;
	signal N3_10_51 : std_logic;
	signal N3_11_52 : std_logic;
	signal N3_12_51 : std_logic;
	signal N3_13_52 : std_logic;
	signal N3_14_51 : std_logic;
	signal N3_15_52 : std_logic;
	signal N3_16_51 : std_logic;
	signal N3_17_52 : std_logic;
	signal N3_18_51 : std_logic;
	signal N3_19_52 : std_logic;
	signal N3_20_51 : std_logic;
	signal N3_21_52 : std_logic;
	signal N3_22_51 : std_logic;
	signal N3_23_52 : std_logic;
	signal N3_0_52 : std_logic;
	signal N3_1_53 : std_logic;
	signal N3_2_52 : std_logic;
	signal N3_3_53 : std_logic;
	signal N3_4_52 : std_logic;
	signal N3_5_53 : std_logic;
	signal N3_6_52 : std_logic;
	signal N3_7_53 : std_logic;
	signal N3_8_52 : std_logic;
	signal N3_9_53 : std_logic;
	signal N3_10_52 : std_logic;
	signal N3_11_53 : std_logic;
	signal N3_12_52 : std_logic;
	signal N3_13_53 : std_logic;
	signal N3_14_52 : std_logic;
	signal N3_15_53 : std_logic;
	signal N3_16_52 : std_logic;
	signal N3_17_53 : std_logic;
	signal N3_18_52 : std_logic;
	signal N3_19_53 : std_logic;
	signal N3_20_52 : std_logic;
	signal N3_21_53 : std_logic;
	signal N3_22_52 : std_logic;
	signal N3_23_53 : std_logic;
	signal N3_0_53 : std_logic;
	signal N3_1_54 : std_logic;
	signal N3_2_53 : std_logic;
	signal N3_3_54 : std_logic;
	signal N3_4_53 : std_logic;
	signal N3_5_54 : std_logic;
	signal N3_6_53 : std_logic;
	signal N3_7_54 : std_logic;
	signal N3_8_53 : std_logic;
	signal N3_9_54 : std_logic;
	signal N3_10_53 : std_logic;
	signal N3_11_54 : std_logic;
	signal N3_12_53 : std_logic;
	signal N3_13_54 : std_logic;
	signal N3_14_53 : std_logic;
	signal N3_15_54 : std_logic;
	signal N3_16_53 : std_logic;
	signal N3_17_54 : std_logic;
	signal N3_18_53 : std_logic;
	signal N3_19_54 : std_logic;
	signal N3_20_53 : std_logic;
	signal N3_21_54 : std_logic;
	signal N3_22_53 : std_logic;
	signal N3_23_54 : std_logic;
	signal N3_0_54 : std_logic;
	signal N3_1_55 : std_logic;
	signal N3_2_54 : std_logic;
	signal N3_3_55 : std_logic;
	signal N3_4_54 : std_logic;
	signal N3_5_55 : std_logic;
	signal N3_6_54 : std_logic;
	signal N3_7_55 : std_logic;
	signal N3_8_54 : std_logic;
	signal N3_9_55 : std_logic;
	signal N3_10_54 : std_logic;
	signal N3_11_55 : std_logic;
	signal N3_12_54 : std_logic;
	signal N3_13_55 : std_logic;
	signal N3_14_54 : std_logic;
	signal N3_15_55 : std_logic;
	signal N3_16_54 : std_logic;
	signal N3_17_55 : std_logic;
	signal N3_18_54 : std_logic;
	signal N3_19_55 : std_logic;
	signal N3_20_54 : std_logic;
	signal N3_21_55 : std_logic;
	signal N3_22_54 : std_logic;
	signal N3_23_55 : std_logic;
	signal N3_0_55 : std_logic;
	signal N3_1_56 : std_logic;
	signal N3_2_55 : std_logic;
	signal N3_3_56 : std_logic;
	signal N3_4_55 : std_logic;
	signal N3_5_56 : std_logic;
	signal N3_6_55 : std_logic;
	signal N3_7_56 : std_logic;
	signal N3_8_55 : std_logic;
	signal N3_9_56 : std_logic;
	signal N3_10_55 : std_logic;
	signal N3_11_56 : std_logic;
	signal N3_12_55 : std_logic;
	signal N3_13_56 : std_logic;
	signal N3_14_55 : std_logic;
	signal N3_15_56 : std_logic;
	signal N3_16_55 : std_logic;
	signal N3_17_56 : std_logic;
	signal N3_18_55 : std_logic;
	signal N3_19_56 : std_logic;
	signal N3_20_55 : std_logic;
	signal N3_21_56 : std_logic;
	signal N3_22_55 : std_logic;
	signal N3_23_56 : std_logic;
	signal N3_0_56 : std_logic;
	signal N3_1_57 : std_logic;
	signal N3_2_56 : std_logic;
	signal N3_3_57 : std_logic;
	signal N3_4_56 : std_logic;
	signal N3_5_57 : std_logic;
	signal N3_6_56 : std_logic;
	signal N3_7_57 : std_logic;
	signal N3_8_56 : std_logic;
	signal N3_9_57 : std_logic;
	signal N3_10_56 : std_logic;
	signal N3_11_57 : std_logic;
	signal N3_12_56 : std_logic;
	signal N3_13_57 : std_logic;
	signal N3_14_56 : std_logic;
	signal N3_15_57 : std_logic;
	signal N3_16_56 : std_logic;
	signal N3_17_57 : std_logic;
	signal N3_18_56 : std_logic;
	signal N3_19_57 : std_logic;
	signal N3_20_56 : std_logic;
	signal N3_21_57 : std_logic;
	signal N3_22_56 : std_logic;
	signal N3_23_57 : std_logic;
	signal N3_0_57 : std_logic;
	signal N3_1_58 : std_logic;
	signal N3_2_57 : std_logic;
	signal N3_3_58 : std_logic;
	signal N3_4_57 : std_logic;
	signal N3_5_58 : std_logic;
	signal N3_6_57 : std_logic;
	signal N3_7_58 : std_logic;
	signal N3_8_57 : std_logic;
	signal N3_9_58 : std_logic;
	signal N3_10_57 : std_logic;
	signal N3_11_58 : std_logic;
	signal N3_12_57 : std_logic;
	signal N3_13_58 : std_logic;
	signal N3_14_57 : std_logic;
	signal N3_15_58 : std_logic;
	signal N3_16_57 : std_logic;
	signal N3_17_58 : std_logic;
	signal N3_18_57 : std_logic;
	signal N3_19_58 : std_logic;
	signal N3_20_57 : std_logic;
	signal N3_21_58 : std_logic;
	signal N3_22_57 : std_logic;
	signal N3_23_58 : std_logic;
	signal N3_0_58 : std_logic;
	signal N3_1_59 : std_logic;
	signal N3_2_58 : std_logic;
	signal N3_3_59 : std_logic;
	signal N3_4_58 : std_logic;
	signal N3_5_59 : std_logic;
	signal N3_6_58 : std_logic;
	signal N3_7_59 : std_logic;
	signal N3_8_58 : std_logic;
	signal N3_9_59 : std_logic;
	signal N3_10_58 : std_logic;
	signal N3_11_59 : std_logic;
	signal N3_12_58 : std_logic;
	signal N3_13_59 : std_logic;
	signal N3_14_58 : std_logic;
	signal N3_15_59 : std_logic;
	signal N3_16_58 : std_logic;
	signal N3_17_59 : std_logic;
	signal N3_18_58 : std_logic;
	signal N3_19_59 : std_logic;
	signal N3_20_58 : std_logic;
	signal N3_21_59 : std_logic;
	signal N3_22_58 : std_logic;
	signal N3_23_59 : std_logic;
	signal N3_0_59 : std_logic;
	signal N3_1_60 : std_logic;
	signal N3_2_59 : std_logic;
	signal N3_3_60 : std_logic;
	signal N3_4_59 : std_logic;
	signal N3_5_60 : std_logic;
	signal N3_6_59 : std_logic;
	signal N3_7_60 : std_logic;
	signal N3_8_59 : std_logic;
	signal N3_9_60 : std_logic;
	signal N3_10_59 : std_logic;
	signal N3_11_60 : std_logic;
	signal N3_12_59 : std_logic;
	signal N3_13_60 : std_logic;
	signal N3_14_59 : std_logic;
	signal N3_15_60 : std_logic;
	signal N3_16_59 : std_logic;
	signal N3_17_60 : std_logic;
	signal N3_18_59 : std_logic;
	signal N3_19_60 : std_logic;
	signal N3_20_59 : std_logic;
	signal N3_21_60 : std_logic;
	signal N3_22_59 : std_logic;
	signal N3_23_60 : std_logic;
	signal N3_0_60 : std_logic;
	signal N3_1_61 : std_logic;
	signal N3_2_60 : std_logic;
	signal N3_3_61 : std_logic;
	signal N3_4_60 : std_logic;
	signal N3_5_61 : std_logic;
	signal N3_6_60 : std_logic;
	signal N3_7_61 : std_logic;
	signal N3_8_60 : std_logic;
	signal N3_9_61 : std_logic;
	signal N3_10_60 : std_logic;
	signal N3_11_61 : std_logic;
	signal N3_12_60 : std_logic;
	signal N3_13_61 : std_logic;
	signal N3_14_60 : std_logic;
	signal N3_15_61 : std_logic;
	signal N3_16_60 : std_logic;
	signal N3_17_61 : std_logic;
	signal N3_18_60 : std_logic;
	signal N3_19_61 : std_logic;
	signal N3_20_60 : std_logic;
	signal N3_21_61 : std_logic;
	signal N3_22_60 : std_logic;
	signal N3_23_61 : std_logic;
	signal N3_0_61 : std_logic;
	signal N3_1_62 : std_logic;
	signal N3_2_61 : std_logic;
	signal N3_3_62 : std_logic;
	signal N3_4_61 : std_logic;
	signal N3_5_62 : std_logic;
	signal N3_6_61 : std_logic;
	signal N3_7_62 : std_logic;
	signal N3_8_61 : std_logic;
	signal N3_9_62 : std_logic;
	signal N3_10_61 : std_logic;
	signal N3_11_62 : std_logic;
	signal N3_12_61 : std_logic;
	signal N3_13_62 : std_logic;
	signal N3_14_61 : std_logic;
	signal N3_15_62 : std_logic;
	signal N3_16_61 : std_logic;
	signal N3_17_62 : std_logic;
	signal N3_18_61 : std_logic;
	signal N3_19_62 : std_logic;
	signal N3_20_61 : std_logic;
	signal N3_21_62 : std_logic;
	signal N3_22_61 : std_logic;
	signal N3_23_62 : std_logic;
	signal N3_0_62 : std_logic;
	signal N3_1_63 : std_logic;
	signal N3_2_62 : std_logic;
	signal N3_3_63 : std_logic;
	signal N3_4_62 : std_logic;
	signal N3_5_63 : std_logic;
	signal N3_6_62 : std_logic;
	signal N3_7_63 : std_logic;
	signal N3_8_62 : std_logic;
	signal N3_9_63 : std_logic;
	signal N3_10_62 : std_logic;
	signal N3_11_63 : std_logic;
	signal N3_12_62 : std_logic;
	signal N3_13_63 : std_logic;
	signal N3_14_62 : std_logic;
	signal N3_15_63 : std_logic;
	signal N3_16_62 : std_logic;
	signal N3_17_63 : std_logic;
	signal N3_18_62 : std_logic;
	signal N3_19_63 : std_logic;
	signal N3_20_62 : std_logic;
	signal N3_21_63 : std_logic;
	signal N3_22_62 : std_logic;
	signal N3_23_63 : std_logic;
	signal N3_0_63 : std_logic;
	signal N3_1_64 : std_logic;
	signal N3_2_63 : std_logic;
	signal N3_3_64 : std_logic;
	signal N3_4_63 : std_logic;
	signal N3_5_64 : std_logic;
	signal N3_6_63 : std_logic;
	signal N3_7_64 : std_logic;
	signal N3_8_63 : std_logic;
	signal N3_9_64 : std_logic;
	signal N3_10_63 : std_logic;
	signal N3_11_64 : std_logic;
	signal N3_12_63 : std_logic;
	signal N3_13_64 : std_logic;
	signal N3_14_63 : std_logic;
	signal N3_15_64 : std_logic;
	signal N3_16_63 : std_logic;
	signal N3_17_64 : std_logic;
	signal N3_18_63 : std_logic;
	signal N3_19_64 : std_logic;
	signal N3_20_63 : std_logic;
	signal N3_21_64 : std_logic;
	signal N3_22_63 : std_logic;
	signal N3_23_64 : std_logic;
	signal N3_0_64 : std_logic;
	signal N3_1_65 : std_logic;
	signal N3_2_64 : std_logic;
	signal N3_3_65 : std_logic;
	signal N3_4_64 : std_logic;
	signal N3_5_65 : std_logic;
	signal N3_6_64 : std_logic;
	signal N3_7_65 : std_logic;
	signal N3_8_64 : std_logic;
	signal N3_9_65 : std_logic;
	signal N3_10_64 : std_logic;
	signal N3_11_65 : std_logic;
	signal N3_12_64 : std_logic;
	signal N3_13_65 : std_logic;
	signal N3_14_64 : std_logic;
	signal N3_15_65 : std_logic;
	signal N3_16_64 : std_logic;
	signal N3_17_65 : std_logic;
	signal N3_18_64 : std_logic;
	signal N3_19_65 : std_logic;
	signal N3_20_64 : std_logic;
	signal N3_21_65 : std_logic;
	signal N3_22_64 : std_logic;
	signal N3_23_65 : std_logic;
	signal N3_0_65 : std_logic;
	signal N3_1_66 : std_logic;
	signal N3_2_65 : std_logic;
	signal N3_3_66 : std_logic;
	signal N3_4_65 : std_logic;
	signal N3_5_66 : std_logic;
	signal N3_6_65 : std_logic;
	signal N3_7_66 : std_logic;
	signal N3_8_65 : std_logic;
	signal N3_9_66 : std_logic;
	signal N3_10_65 : std_logic;
	signal N3_11_66 : std_logic;
	signal N3_12_65 : std_logic;
	signal N3_13_66 : std_logic;
	signal N3_14_65 : std_logic;
	signal N3_15_66 : std_logic;
	signal N3_16_65 : std_logic;
	signal N3_17_66 : std_logic;
	signal N3_18_65 : std_logic;
	signal N3_19_66 : std_logic;
	signal N3_20_65 : std_logic;
	signal N3_21_66 : std_logic;
	signal N3_22_65 : std_logic;
	signal N3_23_66 : std_logic;
	signal N3_0_66 : std_logic;
	signal N3_1_67 : std_logic;
	signal N3_2_66 : std_logic;
	signal N3_3_67 : std_logic;
	signal N3_4_66 : std_logic;
	signal N3_5_67 : std_logic;
	signal N3_6_66 : std_logic;
	signal N3_7_67 : std_logic;
	signal N3_8_66 : std_logic;
	signal N3_9_67 : std_logic;
	signal N3_10_66 : std_logic;
	signal N3_11_67 : std_logic;
	signal N3_12_66 : std_logic;
	signal N3_13_67 : std_logic;
	signal N3_14_66 : std_logic;
	signal N3_15_67 : std_logic;
	signal N3_16_66 : std_logic;
	signal N3_17_67 : std_logic;
	signal N3_18_66 : std_logic;
	signal N3_19_67 : std_logic;
	signal N3_20_66 : std_logic;
	signal N3_21_67 : std_logic;
	signal N3_22_66 : std_logic;
	signal N3_23_67 : std_logic;
	signal N3_0_67 : std_logic;
	signal N3_1_68 : std_logic;
	signal N3_2_67 : std_logic;
	signal N3_3_68 : std_logic;
	signal N3_4_67 : std_logic;
	signal N3_5_68 : std_logic;
	signal N3_6_67 : std_logic;
	signal N3_7_68 : std_logic;
	signal N3_8_67 : std_logic;
	signal N3_9_68 : std_logic;
	signal N3_10_67 : std_logic;
	signal N3_11_68 : std_logic;
	signal N3_12_67 : std_logic;
	signal N3_13_68 : std_logic;
	signal N3_14_67 : std_logic;
	signal N3_15_68 : std_logic;
	signal N3_16_67 : std_logic;
	signal N3_17_68 : std_logic;
	signal N3_18_67 : std_logic;
	signal N3_19_68 : std_logic;
	signal N3_20_67 : std_logic;
	signal N3_21_68 : std_logic;
	signal N3_22_67 : std_logic;
	signal N3_23_68 : std_logic;
	signal N3_0_68 : std_logic;
	signal N3_1_69 : std_logic;
	signal N3_2_68 : std_logic;
	signal N3_3_69 : std_logic;
	signal N3_4_68 : std_logic;
	signal N3_5_69 : std_logic;
	signal N3_6_68 : std_logic;
	signal N3_7_69 : std_logic;
	signal N3_8_68 : std_logic;
	signal N3_9_69 : std_logic;
	signal N3_10_68 : std_logic;
	signal N3_11_69 : std_logic;
	signal N3_12_68 : std_logic;
	signal N3_13_69 : std_logic;
	signal N3_14_68 : std_logic;
	signal N3_15_69 : std_logic;
	signal N3_16_68 : std_logic;
	signal N3_17_69 : std_logic;
	signal N3_18_68 : std_logic;
	signal N3_19_69 : std_logic;
	signal N3_20_68 : std_logic;
	signal N3_21_69 : std_logic;
	signal N3_22_68 : std_logic;
	signal N3_23_69 : std_logic;
	signal N3_0_69 : std_logic;
	signal N3_1_70 : std_logic;
	signal N3_2_69 : std_logic;
	signal N3_3_70 : std_logic;
	signal N3_4_69 : std_logic;
	signal N3_5_70 : std_logic;
	signal N3_6_69 : std_logic;
	signal N3_7_70 : std_logic;
	signal N3_8_69 : std_logic;
	signal N3_9_70 : std_logic;
	signal N3_10_69 : std_logic;
	signal N3_11_70 : std_logic;
	signal N3_12_69 : std_logic;
	signal N3_13_70 : std_logic;
	signal N3_14_69 : std_logic;
	signal N3_15_70 : std_logic;
	signal N3_16_69 : std_logic;
	signal N3_17_70 : std_logic;
	signal N3_18_69 : std_logic;
	signal N3_19_70 : std_logic;
	signal N3_20_69 : std_logic;
	signal N3_21_70 : std_logic;
	signal N3_22_69 : std_logic;
	signal N3_23_70 : std_logic;
	signal N3_0_70 : std_logic;
	signal N3_1_71 : std_logic;
	signal N3_2_70 : std_logic;
	signal N3_3_71 : std_logic;
	signal N3_4_70 : std_logic;
	signal N3_5_71 : std_logic;
	signal N3_6_70 : std_logic;
	signal N3_7_71 : std_logic;
	signal N3_8_70 : std_logic;
	signal N3_9_71 : std_logic;
	signal N3_10_70 : std_logic;
	signal N3_11_71 : std_logic;
	signal N3_12_70 : std_logic;
	signal N3_13_71 : std_logic;
	signal N3_14_70 : std_logic;
	signal N3_15_71 : std_logic;
	signal N3_16_70 : std_logic;
	signal N3_17_71 : std_logic;
	signal N3_18_70 : std_logic;
	signal N3_19_71 : std_logic;
	signal N3_20_70 : std_logic;
	signal N3_21_71 : std_logic;
	signal N3_22_70 : std_logic;
	signal N3_23_71 : std_logic;
	signal N3_0_71 : std_logic;
	signal N3_1_72 : std_logic;
	signal N3_2_71 : std_logic;
	signal N3_3_72 : std_logic;
	signal N3_4_71 : std_logic;
	signal N3_5_72 : std_logic;
	signal N3_6_71 : std_logic;
	signal N3_7_72 : std_logic;
	signal N3_8_71 : std_logic;
	signal N3_9_72 : std_logic;
	signal N3_10_71 : std_logic;
	signal N3_11_72 : std_logic;
	signal N3_12_71 : std_logic;
	signal N3_13_72 : std_logic;
	signal N3_14_71 : std_logic;
	signal N3_15_72 : std_logic;
	signal N3_16_71 : std_logic;
	signal N3_17_72 : std_logic;
	signal N3_18_71 : std_logic;
	signal N3_19_72 : std_logic;
	signal N3_20_71 : std_logic;
	signal N3_21_72 : std_logic;
	signal N3_0_72 : std_logic;
	signal N3_1_73 : std_logic;
	signal N3_2_72 : std_logic;
	signal N3_3_73 : std_logic;
	signal N3_4_72 : std_logic;
	signal N3_5_73 : std_logic;
	signal N3_6_72 : std_logic;
	signal N3_7_73 : std_logic;
	signal N3_8_72 : std_logic;
	signal N3_9_73 : std_logic;
	signal N3_10_72 : std_logic;
	signal N3_11_73 : std_logic;
	signal N3_12_72 : std_logic;
	signal N3_13_73 : std_logic;
	signal N3_14_72 : std_logic;
	signal N3_15_73 : std_logic;
	signal N3_16_72 : std_logic;
	signal N3_17_73 : std_logic;
	signal N3_18_72 : std_logic;
	signal N3_19_73 : std_logic;
	signal N3_0_73 : std_logic;
	signal N3_1_74 : std_logic;
	signal N3_2_73 : std_logic;
	signal N3_3_74 : std_logic;
	signal N3_4_73 : std_logic;
	signal N3_5_74 : std_logic;
	signal N3_6_73 : std_logic;
	signal N3_7_74 : std_logic;
	signal N3_8_73 : std_logic;
	signal N3_9_74 : std_logic;
	signal N3_10_73 : std_logic;
	signal N3_11_74 : std_logic;
	signal N3_12_73 : std_logic;
	signal N3_13_74 : std_logic;
	signal N3_14_73 : std_logic;
	signal N3_15_74 : std_logic;
	signal N3_16_73 : std_logic;
	signal N3_17_74 : std_logic;
	signal N3_0_74 : std_logic;
	signal N3_1_75 : std_logic;
	signal N3_2_74 : std_logic;
	signal N3_3_75 : std_logic;
	signal N3_4_74 : std_logic;
	signal N3_5_75 : std_logic;
	signal N3_6_74 : std_logic;
	signal N3_7_75 : std_logic;
	signal N3_8_74 : std_logic;
	signal N3_9_75 : std_logic;
	signal N3_10_74 : std_logic;
	signal N3_11_75 : std_logic;
	signal N3_12_74 : std_logic;
	signal N3_13_75 : std_logic;
	signal N3_14_74 : std_logic;
	signal N3_15_75 : std_logic;
	signal N3_0_75 : std_logic;
	signal N3_1_76 : std_logic;
	signal N3_2_75 : std_logic;
	signal N3_3_76 : std_logic;
	signal N3_4_75 : std_logic;
	signal N3_5_76 : std_logic;
	signal N3_6_75 : std_logic;
	signal N3_7_76 : std_logic;
	signal N3_8_75 : std_logic;
	signal N3_9_76 : std_logic;
	signal N3_10_75 : std_logic;
	signal N3_11_76 : std_logic;
	signal N3_12_75 : std_logic;
	signal N3_13_76 : std_logic;
	signal N3_0_76 : std_logic;
	signal N3_1_77 : std_logic;
	signal N3_2_76 : std_logic;
	signal N3_3_77 : std_logic;
	signal N3_4_76 : std_logic;
	signal N3_5_77 : std_logic;
	signal N3_6_76 : std_logic;
	signal N3_7_77 : std_logic;
	signal N3_8_76 : std_logic;
	signal N3_9_77 : std_logic;
	signal N3_10_76 : std_logic;
	signal N3_11_77 : std_logic;
	signal N3_0_77 : std_logic;
	signal N3_1_78 : std_logic;
	signal N3_2_77 : std_logic;
	signal N3_3_78 : std_logic;
	signal N3_4_77 : std_logic;
	signal N3_5_78 : std_logic;
	signal N3_6_77 : std_logic;
	signal N3_7_78 : std_logic;
	signal N3_8_77 : std_logic;
	signal N3_9_78 : std_logic;
	signal N3_0_78 : std_logic;
	signal N3_1_79 : std_logic;
	signal N3_2_78 : std_logic;
	signal N3_3_79 : std_logic;
	signal N3_4_78 : std_logic;
	signal N3_5_79 : std_logic;
	signal N3_6_78 : std_logic;
	signal N3_7_79 : std_logic;
	signal N3_0_79 : std_logic;
	signal N3_1_80 : std_logic;
	signal N3_2_79 : std_logic;
	signal N3_3_80 : std_logic;
	signal N3_4_79 : std_logic;
	signal N3_5_80 : std_logic;
	signal N3_0_80 : std_logic;
	signal N3_1_81 : std_logic;
	signal N3_2_80 : std_logic;
	signal N3_3_81 : std_logic;
	signal N3_0_81 : std_logic;
	signal N3_1_82 : std_logic;
	signal N4_0_16 : std_logic;
	signal N4_1_17 : std_logic;
	signal N4_0_17 : std_logic;
	signal N4_1_18 : std_logic;
	signal N4_2_17 : std_logic;
	signal N4_3_18 : std_logic;
	signal N4_0_18 : std_logic;
	signal N4_1_19 : std_logic;
	signal N4_2_18 : std_logic;
	signal N4_3_19 : std_logic;
	signal N4_4_18 : std_logic;
	signal N4_5_19 : std_logic;
	signal N4_0_19 : std_logic;
	signal N4_1_20 : std_logic;
	signal N4_2_19 : std_logic;
	signal N4_3_20 : std_logic;
	signal N4_4_19 : std_logic;
	signal N4_5_20 : std_logic;
	signal N4_6_19 : std_logic;
	signal N4_7_20 : std_logic;
	signal N4_0_20 : std_logic;
	signal N4_1_21 : std_logic;
	signal N4_2_20 : std_logic;
	signal N4_3_21 : std_logic;
	signal N4_4_20 : std_logic;
	signal N4_5_21 : std_logic;
	signal N4_6_20 : std_logic;
	signal N4_7_21 : std_logic;
	signal N4_8_20 : std_logic;
	signal N4_9_21 : std_logic;
	signal N4_0_21 : std_logic;
	signal N4_1_22 : std_logic;
	signal N4_2_21 : std_logic;
	signal N4_3_22 : std_logic;
	signal N4_4_21 : std_logic;
	signal N4_5_22 : std_logic;
	signal N4_6_21 : std_logic;
	signal N4_7_22 : std_logic;
	signal N4_8_21 : std_logic;
	signal N4_9_22 : std_logic;
	signal N4_10_21 : std_logic;
	signal N4_11_22 : std_logic;
	signal N4_0_22 : std_logic;
	signal N4_1_23 : std_logic;
	signal N4_2_22 : std_logic;
	signal N4_3_23 : std_logic;
	signal N4_4_22 : std_logic;
	signal N4_5_23 : std_logic;
	signal N4_6_22 : std_logic;
	signal N4_7_23 : std_logic;
	signal N4_8_22 : std_logic;
	signal N4_9_23 : std_logic;
	signal N4_10_22 : std_logic;
	signal N4_11_23 : std_logic;
	signal N4_12_22 : std_logic;
	signal N4_13_23 : std_logic;
	signal N4_0_23 : std_logic;
	signal N4_1_24 : std_logic;
	signal N4_2_23 : std_logic;
	signal N4_3_24 : std_logic;
	signal N4_4_23 : std_logic;
	signal N4_5_24 : std_logic;
	signal N4_6_23 : std_logic;
	signal N4_7_24 : std_logic;
	signal N4_8_23 : std_logic;
	signal N4_9_24 : std_logic;
	signal N4_10_23 : std_logic;
	signal N4_11_24 : std_logic;
	signal N4_12_23 : std_logic;
	signal N4_13_24 : std_logic;
	signal N4_14_23 : std_logic;
	signal N4_15_24 : std_logic;
	signal N4_0_24 : std_logic;
	signal N4_1_25 : std_logic;
	signal N4_2_24 : std_logic;
	signal N4_3_25 : std_logic;
	signal N4_4_24 : std_logic;
	signal N4_5_25 : std_logic;
	signal N4_6_24 : std_logic;
	signal N4_7_25 : std_logic;
	signal N4_8_24 : std_logic;
	signal N4_9_25 : std_logic;
	signal N4_10_24 : std_logic;
	signal N4_11_25 : std_logic;
	signal N4_12_24 : std_logic;
	signal N4_13_25 : std_logic;
	signal N4_14_24 : std_logic;
	signal N4_15_25 : std_logic;
	signal N4_0_25 : std_logic;
	signal N4_1_26 : std_logic;
	signal N4_2_25 : std_logic;
	signal N4_3_26 : std_logic;
	signal N4_4_25 : std_logic;
	signal N4_5_26 : std_logic;
	signal N4_6_25 : std_logic;
	signal N4_7_26 : std_logic;
	signal N4_8_25 : std_logic;
	signal N4_9_26 : std_logic;
	signal N4_10_25 : std_logic;
	signal N4_11_26 : std_logic;
	signal N4_12_25 : std_logic;
	signal N4_13_26 : std_logic;
	signal N4_14_25 : std_logic;
	signal N4_15_26 : std_logic;
	signal N4_0_26 : std_logic;
	signal N4_1_27 : std_logic;
	signal N4_2_26 : std_logic;
	signal N4_3_27 : std_logic;
	signal N4_4_26 : std_logic;
	signal N4_5_27 : std_logic;
	signal N4_6_26 : std_logic;
	signal N4_7_27 : std_logic;
	signal N4_8_26 : std_logic;
	signal N4_9_27 : std_logic;
	signal N4_10_26 : std_logic;
	signal N4_11_27 : std_logic;
	signal N4_12_26 : std_logic;
	signal N4_13_27 : std_logic;
	signal N4_14_26 : std_logic;
	signal N4_15_27 : std_logic;
	signal N4_0_27 : std_logic;
	signal N4_1_28 : std_logic;
	signal N4_2_27 : std_logic;
	signal N4_3_28 : std_logic;
	signal N4_4_27 : std_logic;
	signal N4_5_28 : std_logic;
	signal N4_6_27 : std_logic;
	signal N4_7_28 : std_logic;
	signal N4_8_27 : std_logic;
	signal N4_9_28 : std_logic;
	signal N4_10_27 : std_logic;
	signal N4_11_28 : std_logic;
	signal N4_12_27 : std_logic;
	signal N4_13_28 : std_logic;
	signal N4_14_27 : std_logic;
	signal N4_15_28 : std_logic;
	signal N4_0_28 : std_logic;
	signal N4_1_29 : std_logic;
	signal N4_2_28 : std_logic;
	signal N4_3_29 : std_logic;
	signal N4_4_28 : std_logic;
	signal N4_5_29 : std_logic;
	signal N4_6_28 : std_logic;
	signal N4_7_29 : std_logic;
	signal N4_8_28 : std_logic;
	signal N4_9_29 : std_logic;
	signal N4_10_28 : std_logic;
	signal N4_11_29 : std_logic;
	signal N4_12_28 : std_logic;
	signal N4_13_29 : std_logic;
	signal N4_14_28 : std_logic;
	signal N4_15_29 : std_logic;
	signal N4_0_29 : std_logic;
	signal N4_1_30 : std_logic;
	signal N4_2_29 : std_logic;
	signal N4_3_30 : std_logic;
	signal N4_4_29 : std_logic;
	signal N4_5_30 : std_logic;
	signal N4_6_29 : std_logic;
	signal N4_7_30 : std_logic;
	signal N4_8_29 : std_logic;
	signal N4_9_30 : std_logic;
	signal N4_10_29 : std_logic;
	signal N4_11_30 : std_logic;
	signal N4_12_29 : std_logic;
	signal N4_13_30 : std_logic;
	signal N4_14_29 : std_logic;
	signal N4_15_30 : std_logic;
	signal N4_0_30 : std_logic;
	signal N4_1_31 : std_logic;
	signal N4_2_30 : std_logic;
	signal N4_3_31 : std_logic;
	signal N4_4_30 : std_logic;
	signal N4_5_31 : std_logic;
	signal N4_6_30 : std_logic;
	signal N4_7_31 : std_logic;
	signal N4_8_30 : std_logic;
	signal N4_9_31 : std_logic;
	signal N4_10_30 : std_logic;
	signal N4_11_31 : std_logic;
	signal N4_12_30 : std_logic;
	signal N4_13_31 : std_logic;
	signal N4_14_30 : std_logic;
	signal N4_15_31 : std_logic;
	signal N4_0_31 : std_logic;
	signal N4_1_32 : std_logic;
	signal N4_2_31 : std_logic;
	signal N4_3_32 : std_logic;
	signal N4_4_31 : std_logic;
	signal N4_5_32 : std_logic;
	signal N4_6_31 : std_logic;
	signal N4_7_32 : std_logic;
	signal N4_8_31 : std_logic;
	signal N4_9_32 : std_logic;
	signal N4_10_31 : std_logic;
	signal N4_11_32 : std_logic;
	signal N4_12_31 : std_logic;
	signal N4_13_32 : std_logic;
	signal N4_14_31 : std_logic;
	signal N4_15_32 : std_logic;
	signal N4_0_32 : std_logic;
	signal N4_1_33 : std_logic;
	signal N4_2_32 : std_logic;
	signal N4_3_33 : std_logic;
	signal N4_4_32 : std_logic;
	signal N4_5_33 : std_logic;
	signal N4_6_32 : std_logic;
	signal N4_7_33 : std_logic;
	signal N4_8_32 : std_logic;
	signal N4_9_33 : std_logic;
	signal N4_10_32 : std_logic;
	signal N4_11_33 : std_logic;
	signal N4_12_32 : std_logic;
	signal N4_13_33 : std_logic;
	signal N4_14_32 : std_logic;
	signal N4_15_33 : std_logic;
	signal N4_0_33 : std_logic;
	signal N4_1_34 : std_logic;
	signal N4_2_33 : std_logic;
	signal N4_3_34 : std_logic;
	signal N4_4_33 : std_logic;
	signal N4_5_34 : std_logic;
	signal N4_6_33 : std_logic;
	signal N4_7_34 : std_logic;
	signal N4_8_33 : std_logic;
	signal N4_9_34 : std_logic;
	signal N4_10_33 : std_logic;
	signal N4_11_34 : std_logic;
	signal N4_12_33 : std_logic;
	signal N4_13_34 : std_logic;
	signal N4_14_33 : std_logic;
	signal N4_15_34 : std_logic;
	signal N4_0_34 : std_logic;
	signal N4_1_35 : std_logic;
	signal N4_2_34 : std_logic;
	signal N4_3_35 : std_logic;
	signal N4_4_34 : std_logic;
	signal N4_5_35 : std_logic;
	signal N4_6_34 : std_logic;
	signal N4_7_35 : std_logic;
	signal N4_8_34 : std_logic;
	signal N4_9_35 : std_logic;
	signal N4_10_34 : std_logic;
	signal N4_11_35 : std_logic;
	signal N4_12_34 : std_logic;
	signal N4_13_35 : std_logic;
	signal N4_14_34 : std_logic;
	signal N4_15_35 : std_logic;
	signal N4_0_35 : std_logic;
	signal N4_1_36 : std_logic;
	signal N4_2_35 : std_logic;
	signal N4_3_36 : std_logic;
	signal N4_4_35 : std_logic;
	signal N4_5_36 : std_logic;
	signal N4_6_35 : std_logic;
	signal N4_7_36 : std_logic;
	signal N4_8_35 : std_logic;
	signal N4_9_36 : std_logic;
	signal N4_10_35 : std_logic;
	signal N4_11_36 : std_logic;
	signal N4_12_35 : std_logic;
	signal N4_13_36 : std_logic;
	signal N4_14_35 : std_logic;
	signal N4_15_36 : std_logic;
	signal N4_0_36 : std_logic;
	signal N4_1_37 : std_logic;
	signal N4_2_36 : std_logic;
	signal N4_3_37 : std_logic;
	signal N4_4_36 : std_logic;
	signal N4_5_37 : std_logic;
	signal N4_6_36 : std_logic;
	signal N4_7_37 : std_logic;
	signal N4_8_36 : std_logic;
	signal N4_9_37 : std_logic;
	signal N4_10_36 : std_logic;
	signal N4_11_37 : std_logic;
	signal N4_12_36 : std_logic;
	signal N4_13_37 : std_logic;
	signal N4_14_36 : std_logic;
	signal N4_15_37 : std_logic;
	signal N4_0_37 : std_logic;
	signal N4_1_38 : std_logic;
	signal N4_2_37 : std_logic;
	signal N4_3_38 : std_logic;
	signal N4_4_37 : std_logic;
	signal N4_5_38 : std_logic;
	signal N4_6_37 : std_logic;
	signal N4_7_38 : std_logic;
	signal N4_8_37 : std_logic;
	signal N4_9_38 : std_logic;
	signal N4_10_37 : std_logic;
	signal N4_11_38 : std_logic;
	signal N4_12_37 : std_logic;
	signal N4_13_38 : std_logic;
	signal N4_14_37 : std_logic;
	signal N4_15_38 : std_logic;
	signal N4_0_38 : std_logic;
	signal N4_1_39 : std_logic;
	signal N4_2_38 : std_logic;
	signal N4_3_39 : std_logic;
	signal N4_4_38 : std_logic;
	signal N4_5_39 : std_logic;
	signal N4_6_38 : std_logic;
	signal N4_7_39 : std_logic;
	signal N4_8_38 : std_logic;
	signal N4_9_39 : std_logic;
	signal N4_10_38 : std_logic;
	signal N4_11_39 : std_logic;
	signal N4_12_38 : std_logic;
	signal N4_13_39 : std_logic;
	signal N4_14_38 : std_logic;
	signal N4_15_39 : std_logic;
	signal N4_0_39 : std_logic;
	signal N4_1_40 : std_logic;
	signal N4_2_39 : std_logic;
	signal N4_3_40 : std_logic;
	signal N4_4_39 : std_logic;
	signal N4_5_40 : std_logic;
	signal N4_6_39 : std_logic;
	signal N4_7_40 : std_logic;
	signal N4_8_39 : std_logic;
	signal N4_9_40 : std_logic;
	signal N4_10_39 : std_logic;
	signal N4_11_40 : std_logic;
	signal N4_12_39 : std_logic;
	signal N4_13_40 : std_logic;
	signal N4_14_39 : std_logic;
	signal N4_15_40 : std_logic;
	signal N4_0_40 : std_logic;
	signal N4_1_41 : std_logic;
	signal N4_2_40 : std_logic;
	signal N4_3_41 : std_logic;
	signal N4_4_40 : std_logic;
	signal N4_5_41 : std_logic;
	signal N4_6_40 : std_logic;
	signal N4_7_41 : std_logic;
	signal N4_8_40 : std_logic;
	signal N4_9_41 : std_logic;
	signal N4_10_40 : std_logic;
	signal N4_11_41 : std_logic;
	signal N4_12_40 : std_logic;
	signal N4_13_41 : std_logic;
	signal N4_14_40 : std_logic;
	signal N4_15_41 : std_logic;
	signal N4_0_41 : std_logic;
	signal N4_1_42 : std_logic;
	signal N4_2_41 : std_logic;
	signal N4_3_42 : std_logic;
	signal N4_4_41 : std_logic;
	signal N4_5_42 : std_logic;
	signal N4_6_41 : std_logic;
	signal N4_7_42 : std_logic;
	signal N4_8_41 : std_logic;
	signal N4_9_42 : std_logic;
	signal N4_10_41 : std_logic;
	signal N4_11_42 : std_logic;
	signal N4_12_41 : std_logic;
	signal N4_13_42 : std_logic;
	signal N4_14_41 : std_logic;
	signal N4_15_42 : std_logic;
	signal N4_0_42 : std_logic;
	signal N4_1_43 : std_logic;
	signal N4_2_42 : std_logic;
	signal N4_3_43 : std_logic;
	signal N4_4_42 : std_logic;
	signal N4_5_43 : std_logic;
	signal N4_6_42 : std_logic;
	signal N4_7_43 : std_logic;
	signal N4_8_42 : std_logic;
	signal N4_9_43 : std_logic;
	signal N4_10_42 : std_logic;
	signal N4_11_43 : std_logic;
	signal N4_12_42 : std_logic;
	signal N4_13_43 : std_logic;
	signal N4_14_42 : std_logic;
	signal N4_15_43 : std_logic;
	signal N4_0_43 : std_logic;
	signal N4_1_44 : std_logic;
	signal N4_2_43 : std_logic;
	signal N4_3_44 : std_logic;
	signal N4_4_43 : std_logic;
	signal N4_5_44 : std_logic;
	signal N4_6_43 : std_logic;
	signal N4_7_44 : std_logic;
	signal N4_8_43 : std_logic;
	signal N4_9_44 : std_logic;
	signal N4_10_43 : std_logic;
	signal N4_11_44 : std_logic;
	signal N4_12_43 : std_logic;
	signal N4_13_44 : std_logic;
	signal N4_14_43 : std_logic;
	signal N4_15_44 : std_logic;
	signal N4_0_44 : std_logic;
	signal N4_1_45 : std_logic;
	signal N4_2_44 : std_logic;
	signal N4_3_45 : std_logic;
	signal N4_4_44 : std_logic;
	signal N4_5_45 : std_logic;
	signal N4_6_44 : std_logic;
	signal N4_7_45 : std_logic;
	signal N4_8_44 : std_logic;
	signal N4_9_45 : std_logic;
	signal N4_10_44 : std_logic;
	signal N4_11_45 : std_logic;
	signal N4_12_44 : std_logic;
	signal N4_13_45 : std_logic;
	signal N4_14_44 : std_logic;
	signal N4_15_45 : std_logic;
	signal N4_0_45 : std_logic;
	signal N4_1_46 : std_logic;
	signal N4_2_45 : std_logic;
	signal N4_3_46 : std_logic;
	signal N4_4_45 : std_logic;
	signal N4_5_46 : std_logic;
	signal N4_6_45 : std_logic;
	signal N4_7_46 : std_logic;
	signal N4_8_45 : std_logic;
	signal N4_9_46 : std_logic;
	signal N4_10_45 : std_logic;
	signal N4_11_46 : std_logic;
	signal N4_12_45 : std_logic;
	signal N4_13_46 : std_logic;
	signal N4_14_45 : std_logic;
	signal N4_15_46 : std_logic;
	signal N4_0_46 : std_logic;
	signal N4_1_47 : std_logic;
	signal N4_2_46 : std_logic;
	signal N4_3_47 : std_logic;
	signal N4_4_46 : std_logic;
	signal N4_5_47 : std_logic;
	signal N4_6_46 : std_logic;
	signal N4_7_47 : std_logic;
	signal N4_8_46 : std_logic;
	signal N4_9_47 : std_logic;
	signal N4_10_46 : std_logic;
	signal N4_11_47 : std_logic;
	signal N4_12_46 : std_logic;
	signal N4_13_47 : std_logic;
	signal N4_14_46 : std_logic;
	signal N4_15_47 : std_logic;
	signal N4_0_47 : std_logic;
	signal N4_1_48 : std_logic;
	signal N4_2_47 : std_logic;
	signal N4_3_48 : std_logic;
	signal N4_4_47 : std_logic;
	signal N4_5_48 : std_logic;
	signal N4_6_47 : std_logic;
	signal N4_7_48 : std_logic;
	signal N4_8_47 : std_logic;
	signal N4_9_48 : std_logic;
	signal N4_10_47 : std_logic;
	signal N4_11_48 : std_logic;
	signal N4_12_47 : std_logic;
	signal N4_13_48 : std_logic;
	signal N4_14_47 : std_logic;
	signal N4_15_48 : std_logic;
	signal N4_0_48 : std_logic;
	signal N4_1_49 : std_logic;
	signal N4_2_48 : std_logic;
	signal N4_3_49 : std_logic;
	signal N4_4_48 : std_logic;
	signal N4_5_49 : std_logic;
	signal N4_6_48 : std_logic;
	signal N4_7_49 : std_logic;
	signal N4_8_48 : std_logic;
	signal N4_9_49 : std_logic;
	signal N4_10_48 : std_logic;
	signal N4_11_49 : std_logic;
	signal N4_12_48 : std_logic;
	signal N4_13_49 : std_logic;
	signal N4_14_48 : std_logic;
	signal N4_15_49 : std_logic;
	signal N4_0_49 : std_logic;
	signal N4_1_50 : std_logic;
	signal N4_2_49 : std_logic;
	signal N4_3_50 : std_logic;
	signal N4_4_49 : std_logic;
	signal N4_5_50 : std_logic;
	signal N4_6_49 : std_logic;
	signal N4_7_50 : std_logic;
	signal N4_8_49 : std_logic;
	signal N4_9_50 : std_logic;
	signal N4_10_49 : std_logic;
	signal N4_11_50 : std_logic;
	signal N4_12_49 : std_logic;
	signal N4_13_50 : std_logic;
	signal N4_14_49 : std_logic;
	signal N4_15_50 : std_logic;
	signal N4_0_50 : std_logic;
	signal N4_1_51 : std_logic;
	signal N4_2_50 : std_logic;
	signal N4_3_51 : std_logic;
	signal N4_4_50 : std_logic;
	signal N4_5_51 : std_logic;
	signal N4_6_50 : std_logic;
	signal N4_7_51 : std_logic;
	signal N4_8_50 : std_logic;
	signal N4_9_51 : std_logic;
	signal N4_10_50 : std_logic;
	signal N4_11_51 : std_logic;
	signal N4_12_50 : std_logic;
	signal N4_13_51 : std_logic;
	signal N4_14_50 : std_logic;
	signal N4_15_51 : std_logic;
	signal N4_0_51 : std_logic;
	signal N4_1_52 : std_logic;
	signal N4_2_51 : std_logic;
	signal N4_3_52 : std_logic;
	signal N4_4_51 : std_logic;
	signal N4_5_52 : std_logic;
	signal N4_6_51 : std_logic;
	signal N4_7_52 : std_logic;
	signal N4_8_51 : std_logic;
	signal N4_9_52 : std_logic;
	signal N4_10_51 : std_logic;
	signal N4_11_52 : std_logic;
	signal N4_12_51 : std_logic;
	signal N4_13_52 : std_logic;
	signal N4_14_51 : std_logic;
	signal N4_15_52 : std_logic;
	signal N4_0_52 : std_logic;
	signal N4_1_53 : std_logic;
	signal N4_2_52 : std_logic;
	signal N4_3_53 : std_logic;
	signal N4_4_52 : std_logic;
	signal N4_5_53 : std_logic;
	signal N4_6_52 : std_logic;
	signal N4_7_53 : std_logic;
	signal N4_8_52 : std_logic;
	signal N4_9_53 : std_logic;
	signal N4_10_52 : std_logic;
	signal N4_11_53 : std_logic;
	signal N4_12_52 : std_logic;
	signal N4_13_53 : std_logic;
	signal N4_14_52 : std_logic;
	signal N4_15_53 : std_logic;
	signal N4_0_53 : std_logic;
	signal N4_1_54 : std_logic;
	signal N4_2_53 : std_logic;
	signal N4_3_54 : std_logic;
	signal N4_4_53 : std_logic;
	signal N4_5_54 : std_logic;
	signal N4_6_53 : std_logic;
	signal N4_7_54 : std_logic;
	signal N4_8_53 : std_logic;
	signal N4_9_54 : std_logic;
	signal N4_10_53 : std_logic;
	signal N4_11_54 : std_logic;
	signal N4_12_53 : std_logic;
	signal N4_13_54 : std_logic;
	signal N4_14_53 : std_logic;
	signal N4_15_54 : std_logic;
	signal N4_0_54 : std_logic;
	signal N4_1_55 : std_logic;
	signal N4_2_54 : std_logic;
	signal N4_3_55 : std_logic;
	signal N4_4_54 : std_logic;
	signal N4_5_55 : std_logic;
	signal N4_6_54 : std_logic;
	signal N4_7_55 : std_logic;
	signal N4_8_54 : std_logic;
	signal N4_9_55 : std_logic;
	signal N4_10_54 : std_logic;
	signal N4_11_55 : std_logic;
	signal N4_12_54 : std_logic;
	signal N4_13_55 : std_logic;
	signal N4_14_54 : std_logic;
	signal N4_15_55 : std_logic;
	signal N4_0_55 : std_logic;
	signal N4_1_56 : std_logic;
	signal N4_2_55 : std_logic;
	signal N4_3_56 : std_logic;
	signal N4_4_55 : std_logic;
	signal N4_5_56 : std_logic;
	signal N4_6_55 : std_logic;
	signal N4_7_56 : std_logic;
	signal N4_8_55 : std_logic;
	signal N4_9_56 : std_logic;
	signal N4_10_55 : std_logic;
	signal N4_11_56 : std_logic;
	signal N4_12_55 : std_logic;
	signal N4_13_56 : std_logic;
	signal N4_14_55 : std_logic;
	signal N4_15_56 : std_logic;
	signal N4_0_56 : std_logic;
	signal N4_1_57 : std_logic;
	signal N4_2_56 : std_logic;
	signal N4_3_57 : std_logic;
	signal N4_4_56 : std_logic;
	signal N4_5_57 : std_logic;
	signal N4_6_56 : std_logic;
	signal N4_7_57 : std_logic;
	signal N4_8_56 : std_logic;
	signal N4_9_57 : std_logic;
	signal N4_10_56 : std_logic;
	signal N4_11_57 : std_logic;
	signal N4_12_56 : std_logic;
	signal N4_13_57 : std_logic;
	signal N4_14_56 : std_logic;
	signal N4_15_57 : std_logic;
	signal N4_0_57 : std_logic;
	signal N4_1_58 : std_logic;
	signal N4_2_57 : std_logic;
	signal N4_3_58 : std_logic;
	signal N4_4_57 : std_logic;
	signal N4_5_58 : std_logic;
	signal N4_6_57 : std_logic;
	signal N4_7_58 : std_logic;
	signal N4_8_57 : std_logic;
	signal N4_9_58 : std_logic;
	signal N4_10_57 : std_logic;
	signal N4_11_58 : std_logic;
	signal N4_12_57 : std_logic;
	signal N4_13_58 : std_logic;
	signal N4_14_57 : std_logic;
	signal N4_15_58 : std_logic;
	signal N4_0_58 : std_logic;
	signal N4_1_59 : std_logic;
	signal N4_2_58 : std_logic;
	signal N4_3_59 : std_logic;
	signal N4_4_58 : std_logic;
	signal N4_5_59 : std_logic;
	signal N4_6_58 : std_logic;
	signal N4_7_59 : std_logic;
	signal N4_8_58 : std_logic;
	signal N4_9_59 : std_logic;
	signal N4_10_58 : std_logic;
	signal N4_11_59 : std_logic;
	signal N4_12_58 : std_logic;
	signal N4_13_59 : std_logic;
	signal N4_14_58 : std_logic;
	signal N4_15_59 : std_logic;
	signal N4_0_59 : std_logic;
	signal N4_1_60 : std_logic;
	signal N4_2_59 : std_logic;
	signal N4_3_60 : std_logic;
	signal N4_4_59 : std_logic;
	signal N4_5_60 : std_logic;
	signal N4_6_59 : std_logic;
	signal N4_7_60 : std_logic;
	signal N4_8_59 : std_logic;
	signal N4_9_60 : std_logic;
	signal N4_10_59 : std_logic;
	signal N4_11_60 : std_logic;
	signal N4_12_59 : std_logic;
	signal N4_13_60 : std_logic;
	signal N4_14_59 : std_logic;
	signal N4_15_60 : std_logic;
	signal N4_0_60 : std_logic;
	signal N4_1_61 : std_logic;
	signal N4_2_60 : std_logic;
	signal N4_3_61 : std_logic;
	signal N4_4_60 : std_logic;
	signal N4_5_61 : std_logic;
	signal N4_6_60 : std_logic;
	signal N4_7_61 : std_logic;
	signal N4_8_60 : std_logic;
	signal N4_9_61 : std_logic;
	signal N4_10_60 : std_logic;
	signal N4_11_61 : std_logic;
	signal N4_12_60 : std_logic;
	signal N4_13_61 : std_logic;
	signal N4_14_60 : std_logic;
	signal N4_15_61 : std_logic;
	signal N4_0_61 : std_logic;
	signal N4_1_62 : std_logic;
	signal N4_2_61 : std_logic;
	signal N4_3_62 : std_logic;
	signal N4_4_61 : std_logic;
	signal N4_5_62 : std_logic;
	signal N4_6_61 : std_logic;
	signal N4_7_62 : std_logic;
	signal N4_8_61 : std_logic;
	signal N4_9_62 : std_logic;
	signal N4_10_61 : std_logic;
	signal N4_11_62 : std_logic;
	signal N4_12_61 : std_logic;
	signal N4_13_62 : std_logic;
	signal N4_14_61 : std_logic;
	signal N4_15_62 : std_logic;
	signal N4_0_62 : std_logic;
	signal N4_1_63 : std_logic;
	signal N4_2_62 : std_logic;
	signal N4_3_63 : std_logic;
	signal N4_4_62 : std_logic;
	signal N4_5_63 : std_logic;
	signal N4_6_62 : std_logic;
	signal N4_7_63 : std_logic;
	signal N4_8_62 : std_logic;
	signal N4_9_63 : std_logic;
	signal N4_10_62 : std_logic;
	signal N4_11_63 : std_logic;
	signal N4_12_62 : std_logic;
	signal N4_13_63 : std_logic;
	signal N4_14_62 : std_logic;
	signal N4_15_63 : std_logic;
	signal N4_0_63 : std_logic;
	signal N4_1_64 : std_logic;
	signal N4_2_63 : std_logic;
	signal N4_3_64 : std_logic;
	signal N4_4_63 : std_logic;
	signal N4_5_64 : std_logic;
	signal N4_6_63 : std_logic;
	signal N4_7_64 : std_logic;
	signal N4_8_63 : std_logic;
	signal N4_9_64 : std_logic;
	signal N4_10_63 : std_logic;
	signal N4_11_64 : std_logic;
	signal N4_12_63 : std_logic;
	signal N4_13_64 : std_logic;
	signal N4_14_63 : std_logic;
	signal N4_15_64 : std_logic;
	signal N4_0_64 : std_logic;
	signal N4_1_65 : std_logic;
	signal N4_2_64 : std_logic;
	signal N4_3_65 : std_logic;
	signal N4_4_64 : std_logic;
	signal N4_5_65 : std_logic;
	signal N4_6_64 : std_logic;
	signal N4_7_65 : std_logic;
	signal N4_8_64 : std_logic;
	signal N4_9_65 : std_logic;
	signal N4_10_64 : std_logic;
	signal N4_11_65 : std_logic;
	signal N4_12_64 : std_logic;
	signal N4_13_65 : std_logic;
	signal N4_14_64 : std_logic;
	signal N4_15_65 : std_logic;
	signal N4_0_65 : std_logic;
	signal N4_1_66 : std_logic;
	signal N4_2_65 : std_logic;
	signal N4_3_66 : std_logic;
	signal N4_4_65 : std_logic;
	signal N4_5_66 : std_logic;
	signal N4_6_65 : std_logic;
	signal N4_7_66 : std_logic;
	signal N4_8_65 : std_logic;
	signal N4_9_66 : std_logic;
	signal N4_10_65 : std_logic;
	signal N4_11_66 : std_logic;
	signal N4_12_65 : std_logic;
	signal N4_13_66 : std_logic;
	signal N4_14_65 : std_logic;
	signal N4_15_66 : std_logic;
	signal N4_0_66 : std_logic;
	signal N4_1_67 : std_logic;
	signal N4_2_66 : std_logic;
	signal N4_3_67 : std_logic;
	signal N4_4_66 : std_logic;
	signal N4_5_67 : std_logic;
	signal N4_6_66 : std_logic;
	signal N4_7_67 : std_logic;
	signal N4_8_66 : std_logic;
	signal N4_9_67 : std_logic;
	signal N4_10_66 : std_logic;
	signal N4_11_67 : std_logic;
	signal N4_12_66 : std_logic;
	signal N4_13_67 : std_logic;
	signal N4_14_66 : std_logic;
	signal N4_15_67 : std_logic;
	signal N4_0_67 : std_logic;
	signal N4_1_68 : std_logic;
	signal N4_2_67 : std_logic;
	signal N4_3_68 : std_logic;
	signal N4_4_67 : std_logic;
	signal N4_5_68 : std_logic;
	signal N4_6_67 : std_logic;
	signal N4_7_68 : std_logic;
	signal N4_8_67 : std_logic;
	signal N4_9_68 : std_logic;
	signal N4_10_67 : std_logic;
	signal N4_11_68 : std_logic;
	signal N4_12_67 : std_logic;
	signal N4_13_68 : std_logic;
	signal N4_14_67 : std_logic;
	signal N4_15_68 : std_logic;
	signal N4_0_68 : std_logic;
	signal N4_1_69 : std_logic;
	signal N4_2_68 : std_logic;
	signal N4_3_69 : std_logic;
	signal N4_4_68 : std_logic;
	signal N4_5_69 : std_logic;
	signal N4_6_68 : std_logic;
	signal N4_7_69 : std_logic;
	signal N4_8_68 : std_logic;
	signal N4_9_69 : std_logic;
	signal N4_10_68 : std_logic;
	signal N4_11_69 : std_logic;
	signal N4_12_68 : std_logic;
	signal N4_13_69 : std_logic;
	signal N4_14_68 : std_logic;
	signal N4_15_69 : std_logic;
	signal N4_0_69 : std_logic;
	signal N4_1_70 : std_logic;
	signal N4_2_69 : std_logic;
	signal N4_3_70 : std_logic;
	signal N4_4_69 : std_logic;
	signal N4_5_70 : std_logic;
	signal N4_6_69 : std_logic;
	signal N4_7_70 : std_logic;
	signal N4_8_69 : std_logic;
	signal N4_9_70 : std_logic;
	signal N4_10_69 : std_logic;
	signal N4_11_70 : std_logic;
	signal N4_12_69 : std_logic;
	signal N4_13_70 : std_logic;
	signal N4_14_69 : std_logic;
	signal N4_15_70 : std_logic;
	signal N4_0_70 : std_logic;
	signal N4_1_71 : std_logic;
	signal N4_2_70 : std_logic;
	signal N4_3_71 : std_logic;
	signal N4_4_70 : std_logic;
	signal N4_5_71 : std_logic;
	signal N4_6_70 : std_logic;
	signal N4_7_71 : std_logic;
	signal N4_8_70 : std_logic;
	signal N4_9_71 : std_logic;
	signal N4_10_70 : std_logic;
	signal N4_11_71 : std_logic;
	signal N4_12_70 : std_logic;
	signal N4_13_71 : std_logic;
	signal N4_14_70 : std_logic;
	signal N4_15_71 : std_logic;
	signal N4_0_71 : std_logic;
	signal N4_1_72 : std_logic;
	signal N4_2_71 : std_logic;
	signal N4_3_72 : std_logic;
	signal N4_4_71 : std_logic;
	signal N4_5_72 : std_logic;
	signal N4_6_71 : std_logic;
	signal N4_7_72 : std_logic;
	signal N4_8_71 : std_logic;
	signal N4_9_72 : std_logic;
	signal N4_10_71 : std_logic;
	signal N4_11_72 : std_logic;
	signal N4_12_71 : std_logic;
	signal N4_13_72 : std_logic;
	signal N4_14_71 : std_logic;
	signal N4_15_72 : std_logic;
	signal N4_0_72 : std_logic;
	signal N4_1_73 : std_logic;
	signal N4_2_72 : std_logic;
	signal N4_3_73 : std_logic;
	signal N4_4_72 : std_logic;
	signal N4_5_73 : std_logic;
	signal N4_6_72 : std_logic;
	signal N4_7_73 : std_logic;
	signal N4_8_72 : std_logic;
	signal N4_9_73 : std_logic;
	signal N4_10_72 : std_logic;
	signal N4_11_73 : std_logic;
	signal N4_12_72 : std_logic;
	signal N4_13_73 : std_logic;
	signal N4_14_72 : std_logic;
	signal N4_15_73 : std_logic;
	signal N4_0_73 : std_logic;
	signal N4_1_74 : std_logic;
	signal N4_2_73 : std_logic;
	signal N4_3_74 : std_logic;
	signal N4_4_73 : std_logic;
	signal N4_5_74 : std_logic;
	signal N4_6_73 : std_logic;
	signal N4_7_74 : std_logic;
	signal N4_8_73 : std_logic;
	signal N4_9_74 : std_logic;
	signal N4_10_73 : std_logic;
	signal N4_11_74 : std_logic;
	signal N4_12_73 : std_logic;
	signal N4_13_74 : std_logic;
	signal N4_14_73 : std_logic;
	signal N4_15_74 : std_logic;
	signal N4_0_74 : std_logic;
	signal N4_1_75 : std_logic;
	signal N4_2_74 : std_logic;
	signal N4_3_75 : std_logic;
	signal N4_4_74 : std_logic;
	signal N4_5_75 : std_logic;
	signal N4_6_74 : std_logic;
	signal N4_7_75 : std_logic;
	signal N4_8_74 : std_logic;
	signal N4_9_75 : std_logic;
	signal N4_10_74 : std_logic;
	signal N4_11_75 : std_logic;
	signal N4_12_74 : std_logic;
	signal N4_13_75 : std_logic;
	signal N4_14_74 : std_logic;
	signal N4_15_75 : std_logic;
	signal N4_0_75 : std_logic;
	signal N4_1_76 : std_logic;
	signal N4_2_75 : std_logic;
	signal N4_3_76 : std_logic;
	signal N4_4_75 : std_logic;
	signal N4_5_76 : std_logic;
	signal N4_6_75 : std_logic;
	signal N4_7_76 : std_logic;
	signal N4_8_75 : std_logic;
	signal N4_9_76 : std_logic;
	signal N4_10_75 : std_logic;
	signal N4_11_76 : std_logic;
	signal N4_12_75 : std_logic;
	signal N4_13_76 : std_logic;
	signal N4_14_75 : std_logic;
	signal N4_15_76 : std_logic;
	signal N4_0_76 : std_logic;
	signal N4_1_77 : std_logic;
	signal N4_2_76 : std_logic;
	signal N4_3_77 : std_logic;
	signal N4_4_76 : std_logic;
	signal N4_5_77 : std_logic;
	signal N4_6_76 : std_logic;
	signal N4_7_77 : std_logic;
	signal N4_8_76 : std_logic;
	signal N4_9_77 : std_logic;
	signal N4_10_76 : std_logic;
	signal N4_11_77 : std_logic;
	signal N4_12_76 : std_logic;
	signal N4_13_77 : std_logic;
	signal N4_14_76 : std_logic;
	signal N4_15_77 : std_logic;
	signal N4_0_77 : std_logic;
	signal N4_1_78 : std_logic;
	signal N4_2_77 : std_logic;
	signal N4_3_78 : std_logic;
	signal N4_4_77 : std_logic;
	signal N4_5_78 : std_logic;
	signal N4_6_77 : std_logic;
	signal N4_7_78 : std_logic;
	signal N4_8_77 : std_logic;
	signal N4_9_78 : std_logic;
	signal N4_10_77 : std_logic;
	signal N4_11_78 : std_logic;
	signal N4_12_77 : std_logic;
	signal N4_13_78 : std_logic;
	signal N4_14_77 : std_logic;
	signal N4_15_78 : std_logic;
	signal N4_0_78 : std_logic;
	signal N4_1_79 : std_logic;
	signal N4_2_78 : std_logic;
	signal N4_3_79 : std_logic;
	signal N4_4_78 : std_logic;
	signal N4_5_79 : std_logic;
	signal N4_6_78 : std_logic;
	signal N4_7_79 : std_logic;
	signal N4_8_78 : std_logic;
	signal N4_9_79 : std_logic;
	signal N4_10_78 : std_logic;
	signal N4_11_79 : std_logic;
	signal N4_12_78 : std_logic;
	signal N4_13_79 : std_logic;
	signal N4_14_78 : std_logic;
	signal N4_15_79 : std_logic;
	signal N4_0_79 : std_logic;
	signal N4_1_80 : std_logic;
	signal N4_2_79 : std_logic;
	signal N4_3_80 : std_logic;
	signal N4_4_79 : std_logic;
	signal N4_5_80 : std_logic;
	signal N4_6_79 : std_logic;
	signal N4_7_80 : std_logic;
	signal N4_8_79 : std_logic;
	signal N4_9_80 : std_logic;
	signal N4_10_79 : std_logic;
	signal N4_11_80 : std_logic;
	signal N4_12_79 : std_logic;
	signal N4_13_80 : std_logic;
	signal N4_14_79 : std_logic;
	signal N4_15_80 : std_logic;
	signal N4_0_80 : std_logic;
	signal N4_1_81 : std_logic;
	signal N4_2_80 : std_logic;
	signal N4_3_81 : std_logic;
	signal N4_4_80 : std_logic;
	signal N4_5_81 : std_logic;
	signal N4_6_80 : std_logic;
	signal N4_7_81 : std_logic;
	signal N4_8_80 : std_logic;
	signal N4_9_81 : std_logic;
	signal N4_10_80 : std_logic;
	signal N4_11_81 : std_logic;
	signal N4_12_80 : std_logic;
	signal N4_13_81 : std_logic;
	signal N4_14_80 : std_logic;
	signal N4_15_81 : std_logic;
	signal N4_0_81 : std_logic;
	signal N4_1_82 : std_logic;
	signal N4_2_81 : std_logic;
	signal N4_3_82 : std_logic;
	signal N4_4_81 : std_logic;
	signal N4_5_82 : std_logic;
	signal N4_6_81 : std_logic;
	signal N4_7_82 : std_logic;
	signal N4_8_81 : std_logic;
	signal N4_9_82 : std_logic;
	signal N4_10_81 : std_logic;
	signal N4_11_82 : std_logic;
	signal N4_12_81 : std_logic;
	signal N4_13_82 : std_logic;
	signal N4_14_81 : std_logic;
	signal N4_15_82 : std_logic;
	signal N4_0_82 : std_logic;
	signal N4_1_83 : std_logic;
	signal N4_2_82 : std_logic;
	signal N4_3_83 : std_logic;
	signal N4_4_82 : std_logic;
	signal N4_5_83 : std_logic;
	signal N4_6_82 : std_logic;
	signal N4_7_83 : std_logic;
	signal N4_8_82 : std_logic;
	signal N4_9_83 : std_logic;
	signal N4_10_82 : std_logic;
	signal N4_11_83 : std_logic;
	signal N4_12_82 : std_logic;
	signal N4_13_83 : std_logic;
	signal N4_14_82 : std_logic;
	signal N4_15_83 : std_logic;
	signal N4_0_83 : std_logic;
	signal N4_1_84 : std_logic;
	signal N4_2_83 : std_logic;
	signal N4_3_84 : std_logic;
	signal N4_4_83 : std_logic;
	signal N4_5_84 : std_logic;
	signal N4_6_83 : std_logic;
	signal N4_7_84 : std_logic;
	signal N4_8_83 : std_logic;
	signal N4_9_84 : std_logic;
	signal N4_10_83 : std_logic;
	signal N4_11_84 : std_logic;
	signal N4_12_83 : std_logic;
	signal N4_13_84 : std_logic;
	signal N4_0_84 : std_logic;
	signal N4_1_85 : std_logic;
	signal N4_2_84 : std_logic;
	signal N4_3_85 : std_logic;
	signal N4_4_84 : std_logic;
	signal N4_5_85 : std_logic;
	signal N4_6_84 : std_logic;
	signal N4_7_85 : std_logic;
	signal N4_8_84 : std_logic;
	signal N4_9_85 : std_logic;
	signal N4_10_84 : std_logic;
	signal N4_11_85 : std_logic;
	signal N4_0_85 : std_logic;
	signal N4_1_86 : std_logic;
	signal N4_2_85 : std_logic;
	signal N4_3_86 : std_logic;
	signal N4_4_85 : std_logic;
	signal N4_5_86 : std_logic;
	signal N4_6_85 : std_logic;
	signal N4_7_86 : std_logic;
	signal N4_8_85 : std_logic;
	signal N4_9_86 : std_logic;
	signal N4_0_86 : std_logic;
	signal N4_1_87 : std_logic;
	signal N4_2_86 : std_logic;
	signal N4_3_87 : std_logic;
	signal N4_4_86 : std_logic;
	signal N4_5_87 : std_logic;
	signal N4_6_86 : std_logic;
	signal N4_7_87 : std_logic;
	signal N4_0_87 : std_logic;
	signal N4_1_88 : std_logic;
	signal N4_2_87 : std_logic;
	signal N4_3_88 : std_logic;
	signal N4_4_87 : std_logic;
	signal N4_5_88 : std_logic;
	signal N4_0_88 : std_logic;
	signal N4_1_89 : std_logic;
	signal N4_2_88 : std_logic;
	signal N4_3_89 : std_logic;
	signal N4_0_89 : std_logic;
	signal N4_1_90 : std_logic;
	signal N5_0_11 : std_logic;
	signal N5_1_12 : std_logic;
	signal N5_0_12 : std_logic;
	signal N5_1_13 : std_logic;
	signal N5_2_12 : std_logic;
	signal N5_3_13 : std_logic;
	signal N5_0_13 : std_logic;
	signal N5_1_14 : std_logic;
	signal N5_2_13 : std_logic;
	signal N5_3_14 : std_logic;
	signal N5_4_13 : std_logic;
	signal N5_5_14 : std_logic;
	signal N5_0_14 : std_logic;
	signal N5_1_15 : std_logic;
	signal N5_2_14 : std_logic;
	signal N5_3_15 : std_logic;
	signal N5_4_14 : std_logic;
	signal N5_5_15 : std_logic;
	signal N5_6_14 : std_logic;
	signal N5_7_15 : std_logic;
	signal N5_0_15 : std_logic;
	signal N5_1_16 : std_logic;
	signal N5_2_15 : std_logic;
	signal N5_3_16 : std_logic;
	signal N5_4_15 : std_logic;
	signal N5_5_16 : std_logic;
	signal N5_6_15 : std_logic;
	signal N5_7_16 : std_logic;
	signal N5_8_15 : std_logic;
	signal N5_9_16 : std_logic;
	signal N5_0_16 : std_logic;
	signal N5_1_17 : std_logic;
	signal N5_2_16 : std_logic;
	signal N5_3_17 : std_logic;
	signal N5_4_16 : std_logic;
	signal N5_5_17 : std_logic;
	signal N5_6_16 : std_logic;
	signal N5_7_17 : std_logic;
	signal N5_8_16 : std_logic;
	signal N5_9_17 : std_logic;
	signal N5_0_17 : std_logic;
	signal N5_1_18 : std_logic;
	signal N5_2_17 : std_logic;
	signal N5_3_18 : std_logic;
	signal N5_4_17 : std_logic;
	signal N5_5_18 : std_logic;
	signal N5_6_17 : std_logic;
	signal N5_7_18 : std_logic;
	signal N5_8_17 : std_logic;
	signal N5_9_18 : std_logic;
	signal N5_0_18 : std_logic;
	signal N5_1_19 : std_logic;
	signal N5_2_18 : std_logic;
	signal N5_3_19 : std_logic;
	signal N5_4_18 : std_logic;
	signal N5_5_19 : std_logic;
	signal N5_6_18 : std_logic;
	signal N5_7_19 : std_logic;
	signal N5_8_18 : std_logic;
	signal N5_9_19 : std_logic;
	signal N5_0_19 : std_logic;
	signal N5_1_20 : std_logic;
	signal N5_2_19 : std_logic;
	signal N5_3_20 : std_logic;
	signal N5_4_19 : std_logic;
	signal N5_5_20 : std_logic;
	signal N5_6_19 : std_logic;
	signal N5_7_20 : std_logic;
	signal N5_8_19 : std_logic;
	signal N5_9_20 : std_logic;
	signal N5_0_20 : std_logic;
	signal N5_1_21 : std_logic;
	signal N5_2_20 : std_logic;
	signal N5_3_21 : std_logic;
	signal N5_4_20 : std_logic;
	signal N5_5_21 : std_logic;
	signal N5_6_20 : std_logic;
	signal N5_7_21 : std_logic;
	signal N5_8_20 : std_logic;
	signal N5_9_21 : std_logic;
	signal N5_0_21 : std_logic;
	signal N5_1_22 : std_logic;
	signal N5_2_21 : std_logic;
	signal N5_3_22 : std_logic;
	signal N5_4_21 : std_logic;
	signal N5_5_22 : std_logic;
	signal N5_6_21 : std_logic;
	signal N5_7_22 : std_logic;
	signal N5_8_21 : std_logic;
	signal N5_9_22 : std_logic;
	signal N5_0_22 : std_logic;
	signal N5_1_23 : std_logic;
	signal N5_2_22 : std_logic;
	signal N5_3_23 : std_logic;
	signal N5_4_22 : std_logic;
	signal N5_5_23 : std_logic;
	signal N5_6_22 : std_logic;
	signal N5_7_23 : std_logic;
	signal N5_8_22 : std_logic;
	signal N5_9_23 : std_logic;
	signal N5_0_23 : std_logic;
	signal N5_1_24 : std_logic;
	signal N5_2_23 : std_logic;
	signal N5_3_24 : std_logic;
	signal N5_4_23 : std_logic;
	signal N5_5_24 : std_logic;
	signal N5_6_23 : std_logic;
	signal N5_7_24 : std_logic;
	signal N5_8_23 : std_logic;
	signal N5_9_24 : std_logic;
	signal N5_0_24 : std_logic;
	signal N5_1_25 : std_logic;
	signal N5_2_24 : std_logic;
	signal N5_3_25 : std_logic;
	signal N5_4_24 : std_logic;
	signal N5_5_25 : std_logic;
	signal N5_6_24 : std_logic;
	signal N5_7_25 : std_logic;
	signal N5_8_24 : std_logic;
	signal N5_9_25 : std_logic;
	signal N5_0_25 : std_logic;
	signal N5_1_26 : std_logic;
	signal N5_2_25 : std_logic;
	signal N5_3_26 : std_logic;
	signal N5_4_25 : std_logic;
	signal N5_5_26 : std_logic;
	signal N5_6_25 : std_logic;
	signal N5_7_26 : std_logic;
	signal N5_8_25 : std_logic;
	signal N5_9_26 : std_logic;
	signal N5_0_26 : std_logic;
	signal N5_1_27 : std_logic;
	signal N5_2_26 : std_logic;
	signal N5_3_27 : std_logic;
	signal N5_4_26 : std_logic;
	signal N5_5_27 : std_logic;
	signal N5_6_26 : std_logic;
	signal N5_7_27 : std_logic;
	signal N5_8_26 : std_logic;
	signal N5_9_27 : std_logic;
	signal N5_0_27 : std_logic;
	signal N5_1_28 : std_logic;
	signal N5_2_27 : std_logic;
	signal N5_3_28 : std_logic;
	signal N5_4_27 : std_logic;
	signal N5_5_28 : std_logic;
	signal N5_6_27 : std_logic;
	signal N5_7_28 : std_logic;
	signal N5_8_27 : std_logic;
	signal N5_9_28 : std_logic;
	signal N5_0_28 : std_logic;
	signal N5_1_29 : std_logic;
	signal N5_2_28 : std_logic;
	signal N5_3_29 : std_logic;
	signal N5_4_28 : std_logic;
	signal N5_5_29 : std_logic;
	signal N5_6_28 : std_logic;
	signal N5_7_29 : std_logic;
	signal N5_8_28 : std_logic;
	signal N5_9_29 : std_logic;
	signal N5_0_29 : std_logic;
	signal N5_1_30 : std_logic;
	signal N5_2_29 : std_logic;
	signal N5_3_30 : std_logic;
	signal N5_4_29 : std_logic;
	signal N5_5_30 : std_logic;
	signal N5_6_29 : std_logic;
	signal N5_7_30 : std_logic;
	signal N5_8_29 : std_logic;
	signal N5_9_30 : std_logic;
	signal N5_0_30 : std_logic;
	signal N5_1_31 : std_logic;
	signal N5_2_30 : std_logic;
	signal N5_3_31 : std_logic;
	signal N5_4_30 : std_logic;
	signal N5_5_31 : std_logic;
	signal N5_6_30 : std_logic;
	signal N5_7_31 : std_logic;
	signal N5_8_30 : std_logic;
	signal N5_9_31 : std_logic;
	signal N5_0_31 : std_logic;
	signal N5_1_32 : std_logic;
	signal N5_2_31 : std_logic;
	signal N5_3_32 : std_logic;
	signal N5_4_31 : std_logic;
	signal N5_5_32 : std_logic;
	signal N5_6_31 : std_logic;
	signal N5_7_32 : std_logic;
	signal N5_8_31 : std_logic;
	signal N5_9_32 : std_logic;
	signal N5_0_32 : std_logic;
	signal N5_1_33 : std_logic;
	signal N5_2_32 : std_logic;
	signal N5_3_33 : std_logic;
	signal N5_4_32 : std_logic;
	signal N5_5_33 : std_logic;
	signal N5_6_32 : std_logic;
	signal N5_7_33 : std_logic;
	signal N5_8_32 : std_logic;
	signal N5_9_33 : std_logic;
	signal N5_0_33 : std_logic;
	signal N5_1_34 : std_logic;
	signal N5_2_33 : std_logic;
	signal N5_3_34 : std_logic;
	signal N5_4_33 : std_logic;
	signal N5_5_34 : std_logic;
	signal N5_6_33 : std_logic;
	signal N5_7_34 : std_logic;
	signal N5_8_33 : std_logic;
	signal N5_9_34 : std_logic;
	signal N5_0_34 : std_logic;
	signal N5_1_35 : std_logic;
	signal N5_2_34 : std_logic;
	signal N5_3_35 : std_logic;
	signal N5_4_34 : std_logic;
	signal N5_5_35 : std_logic;
	signal N5_6_34 : std_logic;
	signal N5_7_35 : std_logic;
	signal N5_8_34 : std_logic;
	signal N5_9_35 : std_logic;
	signal N5_0_35 : std_logic;
	signal N5_1_36 : std_logic;
	signal N5_2_35 : std_logic;
	signal N5_3_36 : std_logic;
	signal N5_4_35 : std_logic;
	signal N5_5_36 : std_logic;
	signal N5_6_35 : std_logic;
	signal N5_7_36 : std_logic;
	signal N5_8_35 : std_logic;
	signal N5_9_36 : std_logic;
	signal N5_0_36 : std_logic;
	signal N5_1_37 : std_logic;
	signal N5_2_36 : std_logic;
	signal N5_3_37 : std_logic;
	signal N5_4_36 : std_logic;
	signal N5_5_37 : std_logic;
	signal N5_6_36 : std_logic;
	signal N5_7_37 : std_logic;
	signal N5_8_36 : std_logic;
	signal N5_9_37 : std_logic;
	signal N5_0_37 : std_logic;
	signal N5_1_38 : std_logic;
	signal N5_2_37 : std_logic;
	signal N5_3_38 : std_logic;
	signal N5_4_37 : std_logic;
	signal N5_5_38 : std_logic;
	signal N5_6_37 : std_logic;
	signal N5_7_38 : std_logic;
	signal N5_8_37 : std_logic;
	signal N5_9_38 : std_logic;
	signal N5_0_38 : std_logic;
	signal N5_1_39 : std_logic;
	signal N5_2_38 : std_logic;
	signal N5_3_39 : std_logic;
	signal N5_4_38 : std_logic;
	signal N5_5_39 : std_logic;
	signal N5_6_38 : std_logic;
	signal N5_7_39 : std_logic;
	signal N5_8_38 : std_logic;
	signal N5_9_39 : std_logic;
	signal N5_0_39 : std_logic;
	signal N5_1_40 : std_logic;
	signal N5_2_39 : std_logic;
	signal N5_3_40 : std_logic;
	signal N5_4_39 : std_logic;
	signal N5_5_40 : std_logic;
	signal N5_6_39 : std_logic;
	signal N5_7_40 : std_logic;
	signal N5_8_39 : std_logic;
	signal N5_9_40 : std_logic;
	signal N5_0_40 : std_logic;
	signal N5_1_41 : std_logic;
	signal N5_2_40 : std_logic;
	signal N5_3_41 : std_logic;
	signal N5_4_40 : std_logic;
	signal N5_5_41 : std_logic;
	signal N5_6_40 : std_logic;
	signal N5_7_41 : std_logic;
	signal N5_8_40 : std_logic;
	signal N5_9_41 : std_logic;
	signal N5_0_41 : std_logic;
	signal N5_1_42 : std_logic;
	signal N5_2_41 : std_logic;
	signal N5_3_42 : std_logic;
	signal N5_4_41 : std_logic;
	signal N5_5_42 : std_logic;
	signal N5_6_41 : std_logic;
	signal N5_7_42 : std_logic;
	signal N5_8_41 : std_logic;
	signal N5_9_42 : std_logic;
	signal N5_0_42 : std_logic;
	signal N5_1_43 : std_logic;
	signal N5_2_42 : std_logic;
	signal N5_3_43 : std_logic;
	signal N5_4_42 : std_logic;
	signal N5_5_43 : std_logic;
	signal N5_6_42 : std_logic;
	signal N5_7_43 : std_logic;
	signal N5_8_42 : std_logic;
	signal N5_9_43 : std_logic;
	signal N5_0_43 : std_logic;
	signal N5_1_44 : std_logic;
	signal N5_2_43 : std_logic;
	signal N5_3_44 : std_logic;
	signal N5_4_43 : std_logic;
	signal N5_5_44 : std_logic;
	signal N5_6_43 : std_logic;
	signal N5_7_44 : std_logic;
	signal N5_8_43 : std_logic;
	signal N5_9_44 : std_logic;
	signal N5_0_44 : std_logic;
	signal N5_1_45 : std_logic;
	signal N5_2_44 : std_logic;
	signal N5_3_45 : std_logic;
	signal N5_4_44 : std_logic;
	signal N5_5_45 : std_logic;
	signal N5_6_44 : std_logic;
	signal N5_7_45 : std_logic;
	signal N5_8_44 : std_logic;
	signal N5_9_45 : std_logic;
	signal N5_0_45 : std_logic;
	signal N5_1_46 : std_logic;
	signal N5_2_45 : std_logic;
	signal N5_3_46 : std_logic;
	signal N5_4_45 : std_logic;
	signal N5_5_46 : std_logic;
	signal N5_6_45 : std_logic;
	signal N5_7_46 : std_logic;
	signal N5_8_45 : std_logic;
	signal N5_9_46 : std_logic;
	signal N5_0_46 : std_logic;
	signal N5_1_47 : std_logic;
	signal N5_2_46 : std_logic;
	signal N5_3_47 : std_logic;
	signal N5_4_46 : std_logic;
	signal N5_5_47 : std_logic;
	signal N5_6_46 : std_logic;
	signal N5_7_47 : std_logic;
	signal N5_8_46 : std_logic;
	signal N5_9_47 : std_logic;
	signal N5_0_47 : std_logic;
	signal N5_1_48 : std_logic;
	signal N5_2_47 : std_logic;
	signal N5_3_48 : std_logic;
	signal N5_4_47 : std_logic;
	signal N5_5_48 : std_logic;
	signal N5_6_47 : std_logic;
	signal N5_7_48 : std_logic;
	signal N5_8_47 : std_logic;
	signal N5_9_48 : std_logic;
	signal N5_0_48 : std_logic;
	signal N5_1_49 : std_logic;
	signal N5_2_48 : std_logic;
	signal N5_3_49 : std_logic;
	signal N5_4_48 : std_logic;
	signal N5_5_49 : std_logic;
	signal N5_6_48 : std_logic;
	signal N5_7_49 : std_logic;
	signal N5_8_48 : std_logic;
	signal N5_9_49 : std_logic;
	signal N5_0_49 : std_logic;
	signal N5_1_50 : std_logic;
	signal N5_2_49 : std_logic;
	signal N5_3_50 : std_logic;
	signal N5_4_49 : std_logic;
	signal N5_5_50 : std_logic;
	signal N5_6_49 : std_logic;
	signal N5_7_50 : std_logic;
	signal N5_8_49 : std_logic;
	signal N5_9_50 : std_logic;
	signal N5_0_50 : std_logic;
	signal N5_1_51 : std_logic;
	signal N5_2_50 : std_logic;
	signal N5_3_51 : std_logic;
	signal N5_4_50 : std_logic;
	signal N5_5_51 : std_logic;
	signal N5_6_50 : std_logic;
	signal N5_7_51 : std_logic;
	signal N5_8_50 : std_logic;
	signal N5_9_51 : std_logic;
	signal N5_0_51 : std_logic;
	signal N5_1_52 : std_logic;
	signal N5_2_51 : std_logic;
	signal N5_3_52 : std_logic;
	signal N5_4_51 : std_logic;
	signal N5_5_52 : std_logic;
	signal N5_6_51 : std_logic;
	signal N5_7_52 : std_logic;
	signal N5_8_51 : std_logic;
	signal N5_9_52 : std_logic;
	signal N5_0_52 : std_logic;
	signal N5_1_53 : std_logic;
	signal N5_2_52 : std_logic;
	signal N5_3_53 : std_logic;
	signal N5_4_52 : std_logic;
	signal N5_5_53 : std_logic;
	signal N5_6_52 : std_logic;
	signal N5_7_53 : std_logic;
	signal N5_8_52 : std_logic;
	signal N5_9_53 : std_logic;
	signal N5_0_53 : std_logic;
	signal N5_1_54 : std_logic;
	signal N5_2_53 : std_logic;
	signal N5_3_54 : std_logic;
	signal N5_4_53 : std_logic;
	signal N5_5_54 : std_logic;
	signal N5_6_53 : std_logic;
	signal N5_7_54 : std_logic;
	signal N5_8_53 : std_logic;
	signal N5_9_54 : std_logic;
	signal N5_0_54 : std_logic;
	signal N5_1_55 : std_logic;
	signal N5_2_54 : std_logic;
	signal N5_3_55 : std_logic;
	signal N5_4_54 : std_logic;
	signal N5_5_55 : std_logic;
	signal N5_6_54 : std_logic;
	signal N5_7_55 : std_logic;
	signal N5_8_54 : std_logic;
	signal N5_9_55 : std_logic;
	signal N5_0_55 : std_logic;
	signal N5_1_56 : std_logic;
	signal N5_2_55 : std_logic;
	signal N5_3_56 : std_logic;
	signal N5_4_55 : std_logic;
	signal N5_5_56 : std_logic;
	signal N5_6_55 : std_logic;
	signal N5_7_56 : std_logic;
	signal N5_8_55 : std_logic;
	signal N5_9_56 : std_logic;
	signal N5_0_56 : std_logic;
	signal N5_1_57 : std_logic;
	signal N5_2_56 : std_logic;
	signal N5_3_57 : std_logic;
	signal N5_4_56 : std_logic;
	signal N5_5_57 : std_logic;
	signal N5_6_56 : std_logic;
	signal N5_7_57 : std_logic;
	signal N5_8_56 : std_logic;
	signal N5_9_57 : std_logic;
	signal N5_0_57 : std_logic;
	signal N5_1_58 : std_logic;
	signal N5_2_57 : std_logic;
	signal N5_3_58 : std_logic;
	signal N5_4_57 : std_logic;
	signal N5_5_58 : std_logic;
	signal N5_6_57 : std_logic;
	signal N5_7_58 : std_logic;
	signal N5_8_57 : std_logic;
	signal N5_9_58 : std_logic;
	signal N5_0_58 : std_logic;
	signal N5_1_59 : std_logic;
	signal N5_2_58 : std_logic;
	signal N5_3_59 : std_logic;
	signal N5_4_58 : std_logic;
	signal N5_5_59 : std_logic;
	signal N5_6_58 : std_logic;
	signal N5_7_59 : std_logic;
	signal N5_8_58 : std_logic;
	signal N5_9_59 : std_logic;
	signal N5_0_59 : std_logic;
	signal N5_1_60 : std_logic;
	signal N5_2_59 : std_logic;
	signal N5_3_60 : std_logic;
	signal N5_4_59 : std_logic;
	signal N5_5_60 : std_logic;
	signal N5_6_59 : std_logic;
	signal N5_7_60 : std_logic;
	signal N5_8_59 : std_logic;
	signal N5_9_60 : std_logic;
	signal N5_0_60 : std_logic;
	signal N5_1_61 : std_logic;
	signal N5_2_60 : std_logic;
	signal N5_3_61 : std_logic;
	signal N5_4_60 : std_logic;
	signal N5_5_61 : std_logic;
	signal N5_6_60 : std_logic;
	signal N5_7_61 : std_logic;
	signal N5_8_60 : std_logic;
	signal N5_9_61 : std_logic;
	signal N5_0_61 : std_logic;
	signal N5_1_62 : std_logic;
	signal N5_2_61 : std_logic;
	signal N5_3_62 : std_logic;
	signal N5_4_61 : std_logic;
	signal N5_5_62 : std_logic;
	signal N5_6_61 : std_logic;
	signal N5_7_62 : std_logic;
	signal N5_8_61 : std_logic;
	signal N5_9_62 : std_logic;
	signal N5_0_62 : std_logic;
	signal N5_1_63 : std_logic;
	signal N5_2_62 : std_logic;
	signal N5_3_63 : std_logic;
	signal N5_4_62 : std_logic;
	signal N5_5_63 : std_logic;
	signal N5_6_62 : std_logic;
	signal N5_7_63 : std_logic;
	signal N5_8_62 : std_logic;
	signal N5_9_63 : std_logic;
	signal N5_0_63 : std_logic;
	signal N5_1_64 : std_logic;
	signal N5_2_63 : std_logic;
	signal N5_3_64 : std_logic;
	signal N5_4_63 : std_logic;
	signal N5_5_64 : std_logic;
	signal N5_6_63 : std_logic;
	signal N5_7_64 : std_logic;
	signal N5_8_63 : std_logic;
	signal N5_9_64 : std_logic;
	signal N5_0_64 : std_logic;
	signal N5_1_65 : std_logic;
	signal N5_2_64 : std_logic;
	signal N5_3_65 : std_logic;
	signal N5_4_64 : std_logic;
	signal N5_5_65 : std_logic;
	signal N5_6_64 : std_logic;
	signal N5_7_65 : std_logic;
	signal N5_8_64 : std_logic;
	signal N5_9_65 : std_logic;
	signal N5_0_65 : std_logic;
	signal N5_1_66 : std_logic;
	signal N5_2_65 : std_logic;
	signal N5_3_66 : std_logic;
	signal N5_4_65 : std_logic;
	signal N5_5_66 : std_logic;
	signal N5_6_65 : std_logic;
	signal N5_7_66 : std_logic;
	signal N5_8_65 : std_logic;
	signal N5_9_66 : std_logic;
	signal N5_0_66 : std_logic;
	signal N5_1_67 : std_logic;
	signal N5_2_66 : std_logic;
	signal N5_3_67 : std_logic;
	signal N5_4_66 : std_logic;
	signal N5_5_67 : std_logic;
	signal N5_6_66 : std_logic;
	signal N5_7_67 : std_logic;
	signal N5_8_66 : std_logic;
	signal N5_9_67 : std_logic;
	signal N5_0_67 : std_logic;
	signal N5_1_68 : std_logic;
	signal N5_2_67 : std_logic;
	signal N5_3_68 : std_logic;
	signal N5_4_67 : std_logic;
	signal N5_5_68 : std_logic;
	signal N5_6_67 : std_logic;
	signal N5_7_68 : std_logic;
	signal N5_8_67 : std_logic;
	signal N5_9_68 : std_logic;
	signal N5_0_68 : std_logic;
	signal N5_1_69 : std_logic;
	signal N5_2_68 : std_logic;
	signal N5_3_69 : std_logic;
	signal N5_4_68 : std_logic;
	signal N5_5_69 : std_logic;
	signal N5_6_68 : std_logic;
	signal N5_7_69 : std_logic;
	signal N5_8_68 : std_logic;
	signal N5_9_69 : std_logic;
	signal N5_0_69 : std_logic;
	signal N5_1_70 : std_logic;
	signal N5_2_69 : std_logic;
	signal N5_3_70 : std_logic;
	signal N5_4_69 : std_logic;
	signal N5_5_70 : std_logic;
	signal N5_6_69 : std_logic;
	signal N5_7_70 : std_logic;
	signal N5_8_69 : std_logic;
	signal N5_9_70 : std_logic;
	signal N5_0_70 : std_logic;
	signal N5_1_71 : std_logic;
	signal N5_2_70 : std_logic;
	signal N5_3_71 : std_logic;
	signal N5_4_70 : std_logic;
	signal N5_5_71 : std_logic;
	signal N5_6_70 : std_logic;
	signal N5_7_71 : std_logic;
	signal N5_8_70 : std_logic;
	signal N5_9_71 : std_logic;
	signal N5_0_71 : std_logic;
	signal N5_1_72 : std_logic;
	signal N5_2_71 : std_logic;
	signal N5_3_72 : std_logic;
	signal N5_4_71 : std_logic;
	signal N5_5_72 : std_logic;
	signal N5_6_71 : std_logic;
	signal N5_7_72 : std_logic;
	signal N5_8_71 : std_logic;
	signal N5_9_72 : std_logic;
	signal N5_0_72 : std_logic;
	signal N5_1_73 : std_logic;
	signal N5_2_72 : std_logic;
	signal N5_3_73 : std_logic;
	signal N5_4_72 : std_logic;
	signal N5_5_73 : std_logic;
	signal N5_6_72 : std_logic;
	signal N5_7_73 : std_logic;
	signal N5_8_72 : std_logic;
	signal N5_9_73 : std_logic;
	signal N5_0_73 : std_logic;
	signal N5_1_74 : std_logic;
	signal N5_2_73 : std_logic;
	signal N5_3_74 : std_logic;
	signal N5_4_73 : std_logic;
	signal N5_5_74 : std_logic;
	signal N5_6_73 : std_logic;
	signal N5_7_74 : std_logic;
	signal N5_8_73 : std_logic;
	signal N5_9_74 : std_logic;
	signal N5_0_74 : std_logic;
	signal N5_1_75 : std_logic;
	signal N5_2_74 : std_logic;
	signal N5_3_75 : std_logic;
	signal N5_4_74 : std_logic;
	signal N5_5_75 : std_logic;
	signal N5_6_74 : std_logic;
	signal N5_7_75 : std_logic;
	signal N5_8_74 : std_logic;
	signal N5_9_75 : std_logic;
	signal N5_0_75 : std_logic;
	signal N5_1_76 : std_logic;
	signal N5_2_75 : std_logic;
	signal N5_3_76 : std_logic;
	signal N5_4_75 : std_logic;
	signal N5_5_76 : std_logic;
	signal N5_6_75 : std_logic;
	signal N5_7_76 : std_logic;
	signal N5_8_75 : std_logic;
	signal N5_9_76 : std_logic;
	signal N5_0_76 : std_logic;
	signal N5_1_77 : std_logic;
	signal N5_2_76 : std_logic;
	signal N5_3_77 : std_logic;
	signal N5_4_76 : std_logic;
	signal N5_5_77 : std_logic;
	signal N5_6_76 : std_logic;
	signal N5_7_77 : std_logic;
	signal N5_8_76 : std_logic;
	signal N5_9_77 : std_logic;
	signal N5_0_77 : std_logic;
	signal N5_1_78 : std_logic;
	signal N5_2_77 : std_logic;
	signal N5_3_78 : std_logic;
	signal N5_4_77 : std_logic;
	signal N5_5_78 : std_logic;
	signal N5_6_77 : std_logic;
	signal N5_7_78 : std_logic;
	signal N5_8_77 : std_logic;
	signal N5_9_78 : std_logic;
	signal N5_0_78 : std_logic;
	signal N5_1_79 : std_logic;
	signal N5_2_78 : std_logic;
	signal N5_3_79 : std_logic;
	signal N5_4_78 : std_logic;
	signal N5_5_79 : std_logic;
	signal N5_6_78 : std_logic;
	signal N5_7_79 : std_logic;
	signal N5_8_78 : std_logic;
	signal N5_9_79 : std_logic;
	signal N5_0_79 : std_logic;
	signal N5_1_80 : std_logic;
	signal N5_2_79 : std_logic;
	signal N5_3_80 : std_logic;
	signal N5_4_79 : std_logic;
	signal N5_5_80 : std_logic;
	signal N5_6_79 : std_logic;
	signal N5_7_80 : std_logic;
	signal N5_8_79 : std_logic;
	signal N5_9_80 : std_logic;
	signal N5_0_80 : std_logic;
	signal N5_1_81 : std_logic;
	signal N5_2_80 : std_logic;
	signal N5_3_81 : std_logic;
	signal N5_4_80 : std_logic;
	signal N5_5_81 : std_logic;
	signal N5_6_80 : std_logic;
	signal N5_7_81 : std_logic;
	signal N5_8_80 : std_logic;
	signal N5_9_81 : std_logic;
	signal N5_0_81 : std_logic;
	signal N5_1_82 : std_logic;
	signal N5_2_81 : std_logic;
	signal N5_3_82 : std_logic;
	signal N5_4_81 : std_logic;
	signal N5_5_82 : std_logic;
	signal N5_6_81 : std_logic;
	signal N5_7_82 : std_logic;
	signal N5_8_81 : std_logic;
	signal N5_9_82 : std_logic;
	signal N5_0_82 : std_logic;
	signal N5_1_83 : std_logic;
	signal N5_2_82 : std_logic;
	signal N5_3_83 : std_logic;
	signal N5_4_82 : std_logic;
	signal N5_5_83 : std_logic;
	signal N5_6_82 : std_logic;
	signal N5_7_83 : std_logic;
	signal N5_8_82 : std_logic;
	signal N5_9_83 : std_logic;
	signal N5_0_83 : std_logic;
	signal N5_1_84 : std_logic;
	signal N5_2_83 : std_logic;
	signal N5_3_84 : std_logic;
	signal N5_4_83 : std_logic;
	signal N5_5_84 : std_logic;
	signal N5_6_83 : std_logic;
	signal N5_7_84 : std_logic;
	signal N5_8_83 : std_logic;
	signal N5_9_84 : std_logic;
	signal N5_0_84 : std_logic;
	signal N5_1_85 : std_logic;
	signal N5_2_84 : std_logic;
	signal N5_3_85 : std_logic;
	signal N5_4_84 : std_logic;
	signal N5_5_85 : std_logic;
	signal N5_6_84 : std_logic;
	signal N5_7_85 : std_logic;
	signal N5_8_84 : std_logic;
	signal N5_9_85 : std_logic;
	signal N5_0_85 : std_logic;
	signal N5_1_86 : std_logic;
	signal N5_2_85 : std_logic;
	signal N5_3_86 : std_logic;
	signal N5_4_85 : std_logic;
	signal N5_5_86 : std_logic;
	signal N5_6_85 : std_logic;
	signal N5_7_86 : std_logic;
	signal N5_8_85 : std_logic;
	signal N5_9_86 : std_logic;
	signal N5_0_86 : std_logic;
	signal N5_1_87 : std_logic;
	signal N5_2_86 : std_logic;
	signal N5_3_87 : std_logic;
	signal N5_4_86 : std_logic;
	signal N5_5_87 : std_logic;
	signal N5_6_86 : std_logic;
	signal N5_7_87 : std_logic;
	signal N5_8_86 : std_logic;
	signal N5_9_87 : std_logic;
	signal N5_0_87 : std_logic;
	signal N5_1_88 : std_logic;
	signal N5_2_87 : std_logic;
	signal N5_3_88 : std_logic;
	signal N5_4_87 : std_logic;
	signal N5_5_88 : std_logic;
	signal N5_6_87 : std_logic;
	signal N5_7_88 : std_logic;
	signal N5_8_87 : std_logic;
	signal N5_9_88 : std_logic;
	signal N5_0_88 : std_logic;
	signal N5_1_89 : std_logic;
	signal N5_2_88 : std_logic;
	signal N5_3_89 : std_logic;
	signal N5_4_88 : std_logic;
	signal N5_5_89 : std_logic;
	signal N5_6_88 : std_logic;
	signal N5_7_89 : std_logic;
	signal N5_8_88 : std_logic;
	signal N5_9_89 : std_logic;
	signal N5_0_89 : std_logic;
	signal N5_1_90 : std_logic;
	signal N5_2_89 : std_logic;
	signal N5_3_90 : std_logic;
	signal N5_4_89 : std_logic;
	signal N5_5_90 : std_logic;
	signal N5_6_89 : std_logic;
	signal N5_7_90 : std_logic;
	signal N5_8_89 : std_logic;
	signal N5_9_90 : std_logic;
	signal N5_0_90 : std_logic;
	signal N5_1_91 : std_logic;
	signal N5_2_90 : std_logic;
	signal N5_3_91 : std_logic;
	signal N5_4_90 : std_logic;
	signal N5_5_91 : std_logic;
	signal N5_6_90 : std_logic;
	signal N5_7_91 : std_logic;
	signal N5_8_90 : std_logic;
	signal N5_9_91 : std_logic;
	signal N5_0_91 : std_logic;
	signal N5_1_92 : std_logic;
	signal N5_2_91 : std_logic;
	signal N5_3_92 : std_logic;
	signal N5_4_91 : std_logic;
	signal N5_5_92 : std_logic;
	signal N5_6_91 : std_logic;
	signal N5_7_92 : std_logic;
	signal N5_0_92 : std_logic;
	signal N5_1_93 : std_logic;
	signal N5_2_92 : std_logic;
	signal N5_3_93 : std_logic;
	signal N5_4_92 : std_logic;
	signal N5_5_93 : std_logic;
	signal N5_0_93 : std_logic;
	signal N5_1_94 : std_logic;
	signal N5_2_93 : std_logic;
	signal N5_3_94 : std_logic;
	signal N5_0_94 : std_logic;
	signal N5_1_95 : std_logic;
	signal N6_0_8 : std_logic;
	signal N6_1_9 : std_logic;
	signal N6_0_9 : std_logic;
	signal N6_1_10 : std_logic;
	signal N6_2_9 : std_logic;
	signal N6_3_10 : std_logic;
	signal N6_0_10 : std_logic;
	signal N6_1_11 : std_logic;
	signal N6_2_10 : std_logic;
	signal N6_3_11 : std_logic;
	signal N6_4_10 : std_logic;
	signal N6_5_11 : std_logic;
	signal N6_0_11 : std_logic;
	signal N6_1_12 : std_logic;
	signal N6_2_11 : std_logic;
	signal N6_3_12 : std_logic;
	signal N6_4_11 : std_logic;
	signal N6_5_12 : std_logic;
	signal N6_0_12 : std_logic;
	signal N6_1_13 : std_logic;
	signal N6_2_12 : std_logic;
	signal N6_3_13 : std_logic;
	signal N6_4_12 : std_logic;
	signal N6_5_13 : std_logic;
	signal N6_0_13 : std_logic;
	signal N6_1_14 : std_logic;
	signal N6_2_13 : std_logic;
	signal N6_3_14 : std_logic;
	signal N6_4_13 : std_logic;
	signal N6_5_14 : std_logic;
	signal N6_0_14 : std_logic;
	signal N6_1_15 : std_logic;
	signal N6_2_14 : std_logic;
	signal N6_3_15 : std_logic;
	signal N6_4_14 : std_logic;
	signal N6_5_15 : std_logic;
	signal N6_0_15 : std_logic;
	signal N6_1_16 : std_logic;
	signal N6_2_15 : std_logic;
	signal N6_3_16 : std_logic;
	signal N6_4_15 : std_logic;
	signal N6_5_16 : std_logic;
	signal N6_0_16 : std_logic;
	signal N6_1_17 : std_logic;
	signal N6_2_16 : std_logic;
	signal N6_3_17 : std_logic;
	signal N6_4_16 : std_logic;
	signal N6_5_17 : std_logic;
	signal N6_0_17 : std_logic;
	signal N6_1_18 : std_logic;
	signal N6_2_17 : std_logic;
	signal N6_3_18 : std_logic;
	signal N6_4_17 : std_logic;
	signal N6_5_18 : std_logic;
	signal N6_0_18 : std_logic;
	signal N6_1_19 : std_logic;
	signal N6_2_18 : std_logic;
	signal N6_3_19 : std_logic;
	signal N6_4_18 : std_logic;
	signal N6_5_19 : std_logic;
	signal N6_0_19 : std_logic;
	signal N6_1_20 : std_logic;
	signal N6_2_19 : std_logic;
	signal N6_3_20 : std_logic;
	signal N6_4_19 : std_logic;
	signal N6_5_20 : std_logic;
	signal N6_0_20 : std_logic;
	signal N6_1_21 : std_logic;
	signal N6_2_20 : std_logic;
	signal N6_3_21 : std_logic;
	signal N6_4_20 : std_logic;
	signal N6_5_21 : std_logic;
	signal N6_0_21 : std_logic;
	signal N6_1_22 : std_logic;
	signal N6_2_21 : std_logic;
	signal N6_3_22 : std_logic;
	signal N6_4_21 : std_logic;
	signal N6_5_22 : std_logic;
	signal N6_0_22 : std_logic;
	signal N6_1_23 : std_logic;
	signal N6_2_22 : std_logic;
	signal N6_3_23 : std_logic;
	signal N6_4_22 : std_logic;
	signal N6_5_23 : std_logic;
	signal N6_0_23 : std_logic;
	signal N6_1_24 : std_logic;
	signal N6_2_23 : std_logic;
	signal N6_3_24 : std_logic;
	signal N6_4_23 : std_logic;
	signal N6_5_24 : std_logic;
	signal N6_0_24 : std_logic;
	signal N6_1_25 : std_logic;
	signal N6_2_24 : std_logic;
	signal N6_3_25 : std_logic;
	signal N6_4_24 : std_logic;
	signal N6_5_25 : std_logic;
	signal N6_0_25 : std_logic;
	signal N6_1_26 : std_logic;
	signal N6_2_25 : std_logic;
	signal N6_3_26 : std_logic;
	signal N6_4_25 : std_logic;
	signal N6_5_26 : std_logic;
	signal N6_0_26 : std_logic;
	signal N6_1_27 : std_logic;
	signal N6_2_26 : std_logic;
	signal N6_3_27 : std_logic;
	signal N6_4_26 : std_logic;
	signal N6_5_27 : std_logic;
	signal N6_0_27 : std_logic;
	signal N6_1_28 : std_logic;
	signal N6_2_27 : std_logic;
	signal N6_3_28 : std_logic;
	signal N6_4_27 : std_logic;
	signal N6_5_28 : std_logic;
	signal N6_0_28 : std_logic;
	signal N6_1_29 : std_logic;
	signal N6_2_28 : std_logic;
	signal N6_3_29 : std_logic;
	signal N6_4_28 : std_logic;
	signal N6_5_29 : std_logic;
	signal N6_0_29 : std_logic;
	signal N6_1_30 : std_logic;
	signal N6_2_29 : std_logic;
	signal N6_3_30 : std_logic;
	signal N6_4_29 : std_logic;
	signal N6_5_30 : std_logic;
	signal N6_0_30 : std_logic;
	signal N6_1_31 : std_logic;
	signal N6_2_30 : std_logic;
	signal N6_3_31 : std_logic;
	signal N6_4_30 : std_logic;
	signal N6_5_31 : std_logic;
	signal N6_0_31 : std_logic;
	signal N6_1_32 : std_logic;
	signal N6_2_31 : std_logic;
	signal N6_3_32 : std_logic;
	signal N6_4_31 : std_logic;
	signal N6_5_32 : std_logic;
	signal N6_0_32 : std_logic;
	signal N6_1_33 : std_logic;
	signal N6_2_32 : std_logic;
	signal N6_3_33 : std_logic;
	signal N6_4_32 : std_logic;
	signal N6_5_33 : std_logic;
	signal N6_0_33 : std_logic;
	signal N6_1_34 : std_logic;
	signal N6_2_33 : std_logic;
	signal N6_3_34 : std_logic;
	signal N6_4_33 : std_logic;
	signal N6_5_34 : std_logic;
	signal N6_0_34 : std_logic;
	signal N6_1_35 : std_logic;
	signal N6_2_34 : std_logic;
	signal N6_3_35 : std_logic;
	signal N6_4_34 : std_logic;
	signal N6_5_35 : std_logic;
	signal N6_0_35 : std_logic;
	signal N6_1_36 : std_logic;
	signal N6_2_35 : std_logic;
	signal N6_3_36 : std_logic;
	signal N6_4_35 : std_logic;
	signal N6_5_36 : std_logic;
	signal N6_0_36 : std_logic;
	signal N6_1_37 : std_logic;
	signal N6_2_36 : std_logic;
	signal N6_3_37 : std_logic;
	signal N6_4_36 : std_logic;
	signal N6_5_37 : std_logic;
	signal N6_0_37 : std_logic;
	signal N6_1_38 : std_logic;
	signal N6_2_37 : std_logic;
	signal N6_3_38 : std_logic;
	signal N6_4_37 : std_logic;
	signal N6_5_38 : std_logic;
	signal N6_0_38 : std_logic;
	signal N6_1_39 : std_logic;
	signal N6_2_38 : std_logic;
	signal N6_3_39 : std_logic;
	signal N6_4_38 : std_logic;
	signal N6_5_39 : std_logic;
	signal N6_0_39 : std_logic;
	signal N6_1_40 : std_logic;
	signal N6_2_39 : std_logic;
	signal N6_3_40 : std_logic;
	signal N6_4_39 : std_logic;
	signal N6_5_40 : std_logic;
	signal N6_0_40 : std_logic;
	signal N6_1_41 : std_logic;
	signal N6_2_40 : std_logic;
	signal N6_3_41 : std_logic;
	signal N6_4_40 : std_logic;
	signal N6_5_41 : std_logic;
	signal N6_0_41 : std_logic;
	signal N6_1_42 : std_logic;
	signal N6_2_41 : std_logic;
	signal N6_3_42 : std_logic;
	signal N6_4_41 : std_logic;
	signal N6_5_42 : std_logic;
	signal N6_0_42 : std_logic;
	signal N6_1_43 : std_logic;
	signal N6_2_42 : std_logic;
	signal N6_3_43 : std_logic;
	signal N6_4_42 : std_logic;
	signal N6_5_43 : std_logic;
	signal N6_0_43 : std_logic;
	signal N6_1_44 : std_logic;
	signal N6_2_43 : std_logic;
	signal N6_3_44 : std_logic;
	signal N6_4_43 : std_logic;
	signal N6_5_44 : std_logic;
	signal N6_0_44 : std_logic;
	signal N6_1_45 : std_logic;
	signal N6_2_44 : std_logic;
	signal N6_3_45 : std_logic;
	signal N6_4_44 : std_logic;
	signal N6_5_45 : std_logic;
	signal N6_0_45 : std_logic;
	signal N6_1_46 : std_logic;
	signal N6_2_45 : std_logic;
	signal N6_3_46 : std_logic;
	signal N6_4_45 : std_logic;
	signal N6_5_46 : std_logic;
	signal N6_0_46 : std_logic;
	signal N6_1_47 : std_logic;
	signal N6_2_46 : std_logic;
	signal N6_3_47 : std_logic;
	signal N6_4_46 : std_logic;
	signal N6_5_47 : std_logic;
	signal N6_0_47 : std_logic;
	signal N6_1_48 : std_logic;
	signal N6_2_47 : std_logic;
	signal N6_3_48 : std_logic;
	signal N6_4_47 : std_logic;
	signal N6_5_48 : std_logic;
	signal N6_0_48 : std_logic;
	signal N6_1_49 : std_logic;
	signal N6_2_48 : std_logic;
	signal N6_3_49 : std_logic;
	signal N6_4_48 : std_logic;
	signal N6_5_49 : std_logic;
	signal N6_0_49 : std_logic;
	signal N6_1_50 : std_logic;
	signal N6_2_49 : std_logic;
	signal N6_3_50 : std_logic;
	signal N6_4_49 : std_logic;
	signal N6_5_50 : std_logic;
	signal N6_0_50 : std_logic;
	signal N6_1_51 : std_logic;
	signal N6_2_50 : std_logic;
	signal N6_3_51 : std_logic;
	signal N6_4_50 : std_logic;
	signal N6_5_51 : std_logic;
	signal N6_0_51 : std_logic;
	signal N6_1_52 : std_logic;
	signal N6_2_51 : std_logic;
	signal N6_3_52 : std_logic;
	signal N6_4_51 : std_logic;
	signal N6_5_52 : std_logic;
	signal N6_0_52 : std_logic;
	signal N6_1_53 : std_logic;
	signal N6_2_52 : std_logic;
	signal N6_3_53 : std_logic;
	signal N6_4_52 : std_logic;
	signal N6_5_53 : std_logic;
	signal N6_0_53 : std_logic;
	signal N6_1_54 : std_logic;
	signal N6_2_53 : std_logic;
	signal N6_3_54 : std_logic;
	signal N6_4_53 : std_logic;
	signal N6_5_54 : std_logic;
	signal N6_0_54 : std_logic;
	signal N6_1_55 : std_logic;
	signal N6_2_54 : std_logic;
	signal N6_3_55 : std_logic;
	signal N6_4_54 : std_logic;
	signal N6_5_55 : std_logic;
	signal N6_0_55 : std_logic;
	signal N6_1_56 : std_logic;
	signal N6_2_55 : std_logic;
	signal N6_3_56 : std_logic;
	signal N6_4_55 : std_logic;
	signal N6_5_56 : std_logic;
	signal N6_0_56 : std_logic;
	signal N6_1_57 : std_logic;
	signal N6_2_56 : std_logic;
	signal N6_3_57 : std_logic;
	signal N6_4_56 : std_logic;
	signal N6_5_57 : std_logic;
	signal N6_0_57 : std_logic;
	signal N6_1_58 : std_logic;
	signal N6_2_57 : std_logic;
	signal N6_3_58 : std_logic;
	signal N6_4_57 : std_logic;
	signal N6_5_58 : std_logic;
	signal N6_0_58 : std_logic;
	signal N6_1_59 : std_logic;
	signal N6_2_58 : std_logic;
	signal N6_3_59 : std_logic;
	signal N6_4_58 : std_logic;
	signal N6_5_59 : std_logic;
	signal N6_0_59 : std_logic;
	signal N6_1_60 : std_logic;
	signal N6_2_59 : std_logic;
	signal N6_3_60 : std_logic;
	signal N6_4_59 : std_logic;
	signal N6_5_60 : std_logic;
	signal N6_0_60 : std_logic;
	signal N6_1_61 : std_logic;
	signal N6_2_60 : std_logic;
	signal N6_3_61 : std_logic;
	signal N6_4_60 : std_logic;
	signal N6_5_61 : std_logic;
	signal N6_0_61 : std_logic;
	signal N6_1_62 : std_logic;
	signal N6_2_61 : std_logic;
	signal N6_3_62 : std_logic;
	signal N6_4_61 : std_logic;
	signal N6_5_62 : std_logic;
	signal N6_0_62 : std_logic;
	signal N6_1_63 : std_logic;
	signal N6_2_62 : std_logic;
	signal N6_3_63 : std_logic;
	signal N6_4_62 : std_logic;
	signal N6_5_63 : std_logic;
	signal N6_0_63 : std_logic;
	signal N6_1_64 : std_logic;
	signal N6_2_63 : std_logic;
	signal N6_3_64 : std_logic;
	signal N6_4_63 : std_logic;
	signal N6_5_64 : std_logic;
	signal N6_0_64 : std_logic;
	signal N6_1_65 : std_logic;
	signal N6_2_64 : std_logic;
	signal N6_3_65 : std_logic;
	signal N6_4_64 : std_logic;
	signal N6_5_65 : std_logic;
	signal N6_0_65 : std_logic;
	signal N6_1_66 : std_logic;
	signal N6_2_65 : std_logic;
	signal N6_3_66 : std_logic;
	signal N6_4_65 : std_logic;
	signal N6_5_66 : std_logic;
	signal N6_0_66 : std_logic;
	signal N6_1_67 : std_logic;
	signal N6_2_66 : std_logic;
	signal N6_3_67 : std_logic;
	signal N6_4_66 : std_logic;
	signal N6_5_67 : std_logic;
	signal N6_0_67 : std_logic;
	signal N6_1_68 : std_logic;
	signal N6_2_67 : std_logic;
	signal N6_3_68 : std_logic;
	signal N6_4_67 : std_logic;
	signal N6_5_68 : std_logic;
	signal N6_0_68 : std_logic;
	signal N6_1_69 : std_logic;
	signal N6_2_68 : std_logic;
	signal N6_3_69 : std_logic;
	signal N6_4_68 : std_logic;
	signal N6_5_69 : std_logic;
	signal N6_0_69 : std_logic;
	signal N6_1_70 : std_logic;
	signal N6_2_69 : std_logic;
	signal N6_3_70 : std_logic;
	signal N6_4_69 : std_logic;
	signal N6_5_70 : std_logic;
	signal N6_0_70 : std_logic;
	signal N6_1_71 : std_logic;
	signal N6_2_70 : std_logic;
	signal N6_3_71 : std_logic;
	signal N6_4_70 : std_logic;
	signal N6_5_71 : std_logic;
	signal N6_0_71 : std_logic;
	signal N6_1_72 : std_logic;
	signal N6_2_71 : std_logic;
	signal N6_3_72 : std_logic;
	signal N6_4_71 : std_logic;
	signal N6_5_72 : std_logic;
	signal N6_0_72 : std_logic;
	signal N6_1_73 : std_logic;
	signal N6_2_72 : std_logic;
	signal N6_3_73 : std_logic;
	signal N6_4_72 : std_logic;
	signal N6_5_73 : std_logic;
	signal N6_0_73 : std_logic;
	signal N6_1_74 : std_logic;
	signal N6_2_73 : std_logic;
	signal N6_3_74 : std_logic;
	signal N6_4_73 : std_logic;
	signal N6_5_74 : std_logic;
	signal N6_0_74 : std_logic;
	signal N6_1_75 : std_logic;
	signal N6_2_74 : std_logic;
	signal N6_3_75 : std_logic;
	signal N6_4_74 : std_logic;
	signal N6_5_75 : std_logic;
	signal N6_0_75 : std_logic;
	signal N6_1_76 : std_logic;
	signal N6_2_75 : std_logic;
	signal N6_3_76 : std_logic;
	signal N6_4_75 : std_logic;
	signal N6_5_76 : std_logic;
	signal N6_0_76 : std_logic;
	signal N6_1_77 : std_logic;
	signal N6_2_76 : std_logic;
	signal N6_3_77 : std_logic;
	signal N6_4_76 : std_logic;
	signal N6_5_77 : std_logic;
	signal N6_0_77 : std_logic;
	signal N6_1_78 : std_logic;
	signal N6_2_77 : std_logic;
	signal N6_3_78 : std_logic;
	signal N6_4_77 : std_logic;
	signal N6_5_78 : std_logic;
	signal N6_0_78 : std_logic;
	signal N6_1_79 : std_logic;
	signal N6_2_78 : std_logic;
	signal N6_3_79 : std_logic;
	signal N6_4_78 : std_logic;
	signal N6_5_79 : std_logic;
	signal N6_0_79 : std_logic;
	signal N6_1_80 : std_logic;
	signal N6_2_79 : std_logic;
	signal N6_3_80 : std_logic;
	signal N6_4_79 : std_logic;
	signal N6_5_80 : std_logic;
	signal N6_0_80 : std_logic;
	signal N6_1_81 : std_logic;
	signal N6_2_80 : std_logic;
	signal N6_3_81 : std_logic;
	signal N6_4_80 : std_logic;
	signal N6_5_81 : std_logic;
	signal N6_0_81 : std_logic;
	signal N6_1_82 : std_logic;
	signal N6_2_81 : std_logic;
	signal N6_3_82 : std_logic;
	signal N6_4_81 : std_logic;
	signal N6_5_82 : std_logic;
	signal N6_0_82 : std_logic;
	signal N6_1_83 : std_logic;
	signal N6_2_82 : std_logic;
	signal N6_3_83 : std_logic;
	signal N6_4_82 : std_logic;
	signal N6_5_83 : std_logic;
	signal N6_0_83 : std_logic;
	signal N6_1_84 : std_logic;
	signal N6_2_83 : std_logic;
	signal N6_3_84 : std_logic;
	signal N6_4_83 : std_logic;
	signal N6_5_84 : std_logic;
	signal N6_0_84 : std_logic;
	signal N6_1_85 : std_logic;
	signal N6_2_84 : std_logic;
	signal N6_3_85 : std_logic;
	signal N6_4_84 : std_logic;
	signal N6_5_85 : std_logic;
	signal N6_0_85 : std_logic;
	signal N6_1_86 : std_logic;
	signal N6_2_85 : std_logic;
	signal N6_3_86 : std_logic;
	signal N6_4_85 : std_logic;
	signal N6_5_86 : std_logic;
	signal N6_0_86 : std_logic;
	signal N6_1_87 : std_logic;
	signal N6_2_86 : std_logic;
	signal N6_3_87 : std_logic;
	signal N6_4_86 : std_logic;
	signal N6_5_87 : std_logic;
	signal N6_0_87 : std_logic;
	signal N6_1_88 : std_logic;
	signal N6_2_87 : std_logic;
	signal N6_3_88 : std_logic;
	signal N6_4_87 : std_logic;
	signal N6_5_88 : std_logic;
	signal N6_0_88 : std_logic;
	signal N6_1_89 : std_logic;
	signal N6_2_88 : std_logic;
	signal N6_3_89 : std_logic;
	signal N6_4_88 : std_logic;
	signal N6_5_89 : std_logic;
	signal N6_0_89 : std_logic;
	signal N6_1_90 : std_logic;
	signal N6_2_89 : std_logic;
	signal N6_3_90 : std_logic;
	signal N6_4_89 : std_logic;
	signal N6_5_90 : std_logic;
	signal N6_0_90 : std_logic;
	signal N6_1_91 : std_logic;
	signal N6_2_90 : std_logic;
	signal N6_3_91 : std_logic;
	signal N6_4_90 : std_logic;
	signal N6_5_91 : std_logic;
	signal N6_0_91 : std_logic;
	signal N6_1_92 : std_logic;
	signal N6_2_91 : std_logic;
	signal N6_3_92 : std_logic;
	signal N6_4_91 : std_logic;
	signal N6_5_92 : std_logic;
	signal N6_0_92 : std_logic;
	signal N6_1_93 : std_logic;
	signal N6_2_92 : std_logic;
	signal N6_3_93 : std_logic;
	signal N6_4_92 : std_logic;
	signal N6_5_93 : std_logic;
	signal N6_0_93 : std_logic;
	signal N6_1_94 : std_logic;
	signal N6_2_93 : std_logic;
	signal N6_3_94 : std_logic;
	signal N6_4_93 : std_logic;
	signal N6_5_94 : std_logic;
	signal N6_0_94 : std_logic;
	signal N6_1_95 : std_logic;
	signal N6_2_94 : std_logic;
	signal N6_3_95 : std_logic;
	signal N6_4_94 : std_logic;
	signal N6_5_95 : std_logic;
	signal N6_0_95 : std_logic;
	signal N6_1_96 : std_logic;
	signal N6_2_95 : std_logic;
	signal N6_3_96 : std_logic;
	signal N6_4_95 : std_logic;
	signal N6_5_96 : std_logic;
	signal N6_0_96 : std_logic;
	signal N6_1_97 : std_logic;
	signal N6_2_96 : std_logic;
	signal N6_3_97 : std_logic;
	signal N6_0_97 : std_logic;
	signal N6_1_98 : std_logic;
	signal N7_0_6 : std_logic;
	signal N7_1_7 : std_logic;
	signal N7_0_7 : std_logic;
	signal N7_1_8 : std_logic;
	signal N7_2_7 : std_logic;
	signal N7_3_8 : std_logic;
	signal N7_0_8 : std_logic;
	signal N7_1_9 : std_logic;
	signal N7_2_8 : std_logic;
	signal N7_3_9 : std_logic;
	signal N7_0_9 : std_logic;
	signal N7_1_10 : std_logic;
	signal N7_2_9 : std_logic;
	signal N7_3_10 : std_logic;
	signal N7_0_10 : std_logic;
	signal N7_1_11 : std_logic;
	signal N7_2_10 : std_logic;
	signal N7_3_11 : std_logic;
	signal N7_0_11 : std_logic;
	signal N7_1_12 : std_logic;
	signal N7_2_11 : std_logic;
	signal N7_3_12 : std_logic;
	signal N7_0_12 : std_logic;
	signal N7_1_13 : std_logic;
	signal N7_2_12 : std_logic;
	signal N7_3_13 : std_logic;
	signal N7_0_13 : std_logic;
	signal N7_1_14 : std_logic;
	signal N7_2_13 : std_logic;
	signal N7_3_14 : std_logic;
	signal N7_0_14 : std_logic;
	signal N7_1_15 : std_logic;
	signal N7_2_14 : std_logic;
	signal N7_3_15 : std_logic;
	signal N7_0_15 : std_logic;
	signal N7_1_16 : std_logic;
	signal N7_2_15 : std_logic;
	signal N7_3_16 : std_logic;
	signal N7_0_16 : std_logic;
	signal N7_1_17 : std_logic;
	signal N7_2_16 : std_logic;
	signal N7_3_17 : std_logic;
	signal N7_0_17 : std_logic;
	signal N7_1_18 : std_logic;
	signal N7_2_17 : std_logic;
	signal N7_3_18 : std_logic;
	signal N7_0_18 : std_logic;
	signal N7_1_19 : std_logic;
	signal N7_2_18 : std_logic;
	signal N7_3_19 : std_logic;
	signal N7_0_19 : std_logic;
	signal N7_1_20 : std_logic;
	signal N7_2_19 : std_logic;
	signal N7_3_20 : std_logic;
	signal N7_0_20 : std_logic;
	signal N7_1_21 : std_logic;
	signal N7_2_20 : std_logic;
	signal N7_3_21 : std_logic;
	signal N7_0_21 : std_logic;
	signal N7_1_22 : std_logic;
	signal N7_2_21 : std_logic;
	signal N7_3_22 : std_logic;
	signal N7_0_22 : std_logic;
	signal N7_1_23 : std_logic;
	signal N7_2_22 : std_logic;
	signal N7_3_23 : std_logic;
	signal N7_0_23 : std_logic;
	signal N7_1_24 : std_logic;
	signal N7_2_23 : std_logic;
	signal N7_3_24 : std_logic;
	signal N7_0_24 : std_logic;
	signal N7_1_25 : std_logic;
	signal N7_2_24 : std_logic;
	signal N7_3_25 : std_logic;
	signal N7_0_25 : std_logic;
	signal N7_1_26 : std_logic;
	signal N7_2_25 : std_logic;
	signal N7_3_26 : std_logic;
	signal N7_0_26 : std_logic;
	signal N7_1_27 : std_logic;
	signal N7_2_26 : std_logic;
	signal N7_3_27 : std_logic;
	signal N7_0_27 : std_logic;
	signal N7_1_28 : std_logic;
	signal N7_2_27 : std_logic;
	signal N7_3_28 : std_logic;
	signal N7_0_28 : std_logic;
	signal N7_1_29 : std_logic;
	signal N7_2_28 : std_logic;
	signal N7_3_29 : std_logic;
	signal N7_0_29 : std_logic;
	signal N7_1_30 : std_logic;
	signal N7_2_29 : std_logic;
	signal N7_3_30 : std_logic;
	signal N7_0_30 : std_logic;
	signal N7_1_31 : std_logic;
	signal N7_2_30 : std_logic;
	signal N7_3_31 : std_logic;
	signal N7_0_31 : std_logic;
	signal N7_1_32 : std_logic;
	signal N7_2_31 : std_logic;
	signal N7_3_32 : std_logic;
	signal N7_0_32 : std_logic;
	signal N7_1_33 : std_logic;
	signal N7_2_32 : std_logic;
	signal N7_3_33 : std_logic;
	signal N7_0_33 : std_logic;
	signal N7_1_34 : std_logic;
	signal N7_2_33 : std_logic;
	signal N7_3_34 : std_logic;
	signal N7_0_34 : std_logic;
	signal N7_1_35 : std_logic;
	signal N7_2_34 : std_logic;
	signal N7_3_35 : std_logic;
	signal N7_0_35 : std_logic;
	signal N7_1_36 : std_logic;
	signal N7_2_35 : std_logic;
	signal N7_3_36 : std_logic;
	signal N7_0_36 : std_logic;
	signal N7_1_37 : std_logic;
	signal N7_2_36 : std_logic;
	signal N7_3_37 : std_logic;
	signal N7_0_37 : std_logic;
	signal N7_1_38 : std_logic;
	signal N7_2_37 : std_logic;
	signal N7_3_38 : std_logic;
	signal N7_0_38 : std_logic;
	signal N7_1_39 : std_logic;
	signal N7_2_38 : std_logic;
	signal N7_3_39 : std_logic;
	signal N7_0_39 : std_logic;
	signal N7_1_40 : std_logic;
	signal N7_2_39 : std_logic;
	signal N7_3_40 : std_logic;
	signal N7_0_40 : std_logic;
	signal N7_1_41 : std_logic;
	signal N7_2_40 : std_logic;
	signal N7_3_41 : std_logic;
	signal N7_0_41 : std_logic;
	signal N7_1_42 : std_logic;
	signal N7_2_41 : std_logic;
	signal N7_3_42 : std_logic;
	signal N7_0_42 : std_logic;
	signal N7_1_43 : std_logic;
	signal N7_2_42 : std_logic;
	signal N7_3_43 : std_logic;
	signal N7_0_43 : std_logic;
	signal N7_1_44 : std_logic;
	signal N7_2_43 : std_logic;
	signal N7_3_44 : std_logic;
	signal N7_0_44 : std_logic;
	signal N7_1_45 : std_logic;
	signal N7_2_44 : std_logic;
	signal N7_3_45 : std_logic;
	signal N7_0_45 : std_logic;
	signal N7_1_46 : std_logic;
	signal N7_2_45 : std_logic;
	signal N7_3_46 : std_logic;
	signal N7_0_46 : std_logic;
	signal N7_1_47 : std_logic;
	signal N7_2_46 : std_logic;
	signal N7_3_47 : std_logic;
	signal N7_0_47 : std_logic;
	signal N7_1_48 : std_logic;
	signal N7_2_47 : std_logic;
	signal N7_3_48 : std_logic;
	signal N7_0_48 : std_logic;
	signal N7_1_49 : std_logic;
	signal N7_2_48 : std_logic;
	signal N7_3_49 : std_logic;
	signal N7_0_49 : std_logic;
	signal N7_1_50 : std_logic;
	signal N7_2_49 : std_logic;
	signal N7_3_50 : std_logic;
	signal N7_0_50 : std_logic;
	signal N7_1_51 : std_logic;
	signal N7_2_50 : std_logic;
	signal N7_3_51 : std_logic;
	signal N7_0_51 : std_logic;
	signal N7_1_52 : std_logic;
	signal N7_2_51 : std_logic;
	signal N7_3_52 : std_logic;
	signal N7_0_52 : std_logic;
	signal N7_1_53 : std_logic;
	signal N7_2_52 : std_logic;
	signal N7_3_53 : std_logic;
	signal N7_0_53 : std_logic;
	signal N7_1_54 : std_logic;
	signal N7_2_53 : std_logic;
	signal N7_3_54 : std_logic;
	signal N7_0_54 : std_logic;
	signal N7_1_55 : std_logic;
	signal N7_2_54 : std_logic;
	signal N7_3_55 : std_logic;
	signal N7_0_55 : std_logic;
	signal N7_1_56 : std_logic;
	signal N7_2_55 : std_logic;
	signal N7_3_56 : std_logic;
	signal N7_0_56 : std_logic;
	signal N7_1_57 : std_logic;
	signal N7_2_56 : std_logic;
	signal N7_3_57 : std_logic;
	signal N7_0_57 : std_logic;
	signal N7_1_58 : std_logic;
	signal N7_2_57 : std_logic;
	signal N7_3_58 : std_logic;
	signal N7_0_58 : std_logic;
	signal N7_1_59 : std_logic;
	signal N7_2_58 : std_logic;
	signal N7_3_59 : std_logic;
	signal N7_0_59 : std_logic;
	signal N7_1_60 : std_logic;
	signal N7_2_59 : std_logic;
	signal N7_3_60 : std_logic;
	signal N7_0_60 : std_logic;
	signal N7_1_61 : std_logic;
	signal N7_2_60 : std_logic;
	signal N7_3_61 : std_logic;
	signal N7_0_61 : std_logic;
	signal N7_1_62 : std_logic;
	signal N7_2_61 : std_logic;
	signal N7_3_62 : std_logic;
	signal N7_0_62 : std_logic;
	signal N7_1_63 : std_logic;
	signal N7_2_62 : std_logic;
	signal N7_3_63 : std_logic;
	signal N7_0_63 : std_logic;
	signal N7_1_64 : std_logic;
	signal N7_2_63 : std_logic;
	signal N7_3_64 : std_logic;
	signal N7_0_64 : std_logic;
	signal N7_1_65 : std_logic;
	signal N7_2_64 : std_logic;
	signal N7_3_65 : std_logic;
	signal N7_0_65 : std_logic;
	signal N7_1_66 : std_logic;
	signal N7_2_65 : std_logic;
	signal N7_3_66 : std_logic;
	signal N7_0_66 : std_logic;
	signal N7_1_67 : std_logic;
	signal N7_2_66 : std_logic;
	signal N7_3_67 : std_logic;
	signal N7_0_67 : std_logic;
	signal N7_1_68 : std_logic;
	signal N7_2_67 : std_logic;
	signal N7_3_68 : std_logic;
	signal N7_0_68 : std_logic;
	signal N7_1_69 : std_logic;
	signal N7_2_68 : std_logic;
	signal N7_3_69 : std_logic;
	signal N7_0_69 : std_logic;
	signal N7_1_70 : std_logic;
	signal N7_2_69 : std_logic;
	signal N7_3_70 : std_logic;
	signal N7_0_70 : std_logic;
	signal N7_1_71 : std_logic;
	signal N7_2_70 : std_logic;
	signal N7_3_71 : std_logic;
	signal N7_0_71 : std_logic;
	signal N7_1_72 : std_logic;
	signal N7_2_71 : std_logic;
	signal N7_3_72 : std_logic;
	signal N7_0_72 : std_logic;
	signal N7_1_73 : std_logic;
	signal N7_2_72 : std_logic;
	signal N7_3_73 : std_logic;
	signal N7_0_73 : std_logic;
	signal N7_1_74 : std_logic;
	signal N7_2_73 : std_logic;
	signal N7_3_74 : std_logic;
	signal N7_0_74 : std_logic;
	signal N7_1_75 : std_logic;
	signal N7_2_74 : std_logic;
	signal N7_3_75 : std_logic;
	signal N7_0_75 : std_logic;
	signal N7_1_76 : std_logic;
	signal N7_2_75 : std_logic;
	signal N7_3_76 : std_logic;
	signal N7_0_76 : std_logic;
	signal N7_1_77 : std_logic;
	signal N7_2_76 : std_logic;
	signal N7_3_77 : std_logic;
	signal N7_0_77 : std_logic;
	signal N7_1_78 : std_logic;
	signal N7_2_77 : std_logic;
	signal N7_3_78 : std_logic;
	signal N7_0_78 : std_logic;
	signal N7_1_79 : std_logic;
	signal N7_2_78 : std_logic;
	signal N7_3_79 : std_logic;
	signal N7_0_79 : std_logic;
	signal N7_1_80 : std_logic;
	signal N7_2_79 : std_logic;
	signal N7_3_80 : std_logic;
	signal N7_0_80 : std_logic;
	signal N7_1_81 : std_logic;
	signal N7_2_80 : std_logic;
	signal N7_3_81 : std_logic;
	signal N7_0_81 : std_logic;
	signal N7_1_82 : std_logic;
	signal N7_2_81 : std_logic;
	signal N7_3_82 : std_logic;
	signal N7_0_82 : std_logic;
	signal N7_1_83 : std_logic;
	signal N7_2_82 : std_logic;
	signal N7_3_83 : std_logic;
	signal N7_0_83 : std_logic;
	signal N7_1_84 : std_logic;
	signal N7_2_83 : std_logic;
	signal N7_3_84 : std_logic;
	signal N7_0_84 : std_logic;
	signal N7_1_85 : std_logic;
	signal N7_2_84 : std_logic;
	signal N7_3_85 : std_logic;
	signal N7_0_85 : std_logic;
	signal N7_1_86 : std_logic;
	signal N7_2_85 : std_logic;
	signal N7_3_86 : std_logic;
	signal N7_0_86 : std_logic;
	signal N7_1_87 : std_logic;
	signal N7_2_86 : std_logic;
	signal N7_3_87 : std_logic;
	signal N7_0_87 : std_logic;
	signal N7_1_88 : std_logic;
	signal N7_2_87 : std_logic;
	signal N7_3_88 : std_logic;
	signal N7_0_88 : std_logic;
	signal N7_1_89 : std_logic;
	signal N7_2_88 : std_logic;
	signal N7_3_89 : std_logic;
	signal N7_0_89 : std_logic;
	signal N7_1_90 : std_logic;
	signal N7_2_89 : std_logic;
	signal N7_3_90 : std_logic;
	signal N7_0_90 : std_logic;
	signal N7_1_91 : std_logic;
	signal N7_2_90 : std_logic;
	signal N7_3_91 : std_logic;
	signal N7_0_91 : std_logic;
	signal N7_1_92 : std_logic;
	signal N7_2_91 : std_logic;
	signal N7_3_92 : std_logic;
	signal N7_0_92 : std_logic;
	signal N7_1_93 : std_logic;
	signal N7_2_92 : std_logic;
	signal N7_3_93 : std_logic;
	signal N7_0_93 : std_logic;
	signal N7_1_94 : std_logic;
	signal N7_2_93 : std_logic;
	signal N7_3_94 : std_logic;
	signal N7_0_94 : std_logic;
	signal N7_1_95 : std_logic;
	signal N7_2_94 : std_logic;
	signal N7_3_95 : std_logic;
	signal N7_0_95 : std_logic;
	signal N7_1_96 : std_logic;
	signal N7_2_95 : std_logic;
	signal N7_3_96 : std_logic;
	signal N7_0_96 : std_logic;
	signal N7_1_97 : std_logic;
	signal N7_2_96 : std_logic;
	signal N7_3_97 : std_logic;
	signal N7_0_97 : std_logic;
	signal N7_1_98 : std_logic;
	signal N7_2_97 : std_logic;
	signal N7_3_98 : std_logic;
	signal N7_0_98 : std_logic;
	signal N7_1_99 : std_logic;
	signal N7_2_98 : std_logic;
	signal N7_3_99 : std_logic;
	signal N7_0_99 : std_logic;
	signal N7_1_100 : std_logic;
	signal N8_0_4 : std_logic;
	signal N8_1_5 : std_logic;
	signal N8_0_5 : std_logic;
	signal N8_1_6 : std_logic;
	signal N8_2_5 : std_logic;
	signal N8_3_6 : std_logic;
	signal N8_0_6 : std_logic;
	signal N8_1_7 : std_logic;
	signal N8_2_6 : std_logic;
	signal N8_3_7 : std_logic;
	signal N8_0_7 : std_logic;
	signal N8_1_8 : std_logic;
	signal N8_2_7 : std_logic;
	signal N8_3_8 : std_logic;
	signal N8_0_8 : std_logic;
	signal N8_1_9 : std_logic;
	signal N8_2_8 : std_logic;
	signal N8_3_9 : std_logic;
	signal N8_0_9 : std_logic;
	signal N8_1_10 : std_logic;
	signal N8_2_9 : std_logic;
	signal N8_3_10 : std_logic;
	signal N8_0_10 : std_logic;
	signal N8_1_11 : std_logic;
	signal N8_2_10 : std_logic;
	signal N8_3_11 : std_logic;
	signal N8_0_11 : std_logic;
	signal N8_1_12 : std_logic;
	signal N8_2_11 : std_logic;
	signal N8_3_12 : std_logic;
	signal N8_0_12 : std_logic;
	signal N8_1_13 : std_logic;
	signal N8_2_12 : std_logic;
	signal N8_3_13 : std_logic;
	signal N8_0_13 : std_logic;
	signal N8_1_14 : std_logic;
	signal N8_2_13 : std_logic;
	signal N8_3_14 : std_logic;
	signal N8_0_14 : std_logic;
	signal N8_1_15 : std_logic;
	signal N8_2_14 : std_logic;
	signal N8_3_15 : std_logic;
	signal N8_0_15 : std_logic;
	signal N8_1_16 : std_logic;
	signal N8_2_15 : std_logic;
	signal N8_3_16 : std_logic;
	signal N8_0_16 : std_logic;
	signal N8_1_17 : std_logic;
	signal N8_2_16 : std_logic;
	signal N8_3_17 : std_logic;
	signal N8_0_17 : std_logic;
	signal N8_1_18 : std_logic;
	signal N8_2_17 : std_logic;
	signal N8_3_18 : std_logic;
	signal N8_0_18 : std_logic;
	signal N8_1_19 : std_logic;
	signal N8_2_18 : std_logic;
	signal N8_3_19 : std_logic;
	signal N8_0_19 : std_logic;
	signal N8_1_20 : std_logic;
	signal N8_2_19 : std_logic;
	signal N8_3_20 : std_logic;
	signal N8_0_20 : std_logic;
	signal N8_1_21 : std_logic;
	signal N8_2_20 : std_logic;
	signal N8_3_21 : std_logic;
	signal N8_0_21 : std_logic;
	signal N8_1_22 : std_logic;
	signal N8_2_21 : std_logic;
	signal N8_3_22 : std_logic;
	signal N8_0_22 : std_logic;
	signal N8_1_23 : std_logic;
	signal N8_2_22 : std_logic;
	signal N8_3_23 : std_logic;
	signal N8_0_23 : std_logic;
	signal N8_1_24 : std_logic;
	signal N8_2_23 : std_logic;
	signal N8_3_24 : std_logic;
	signal N8_0_24 : std_logic;
	signal N8_1_25 : std_logic;
	signal N8_2_24 : std_logic;
	signal N8_3_25 : std_logic;
	signal N8_0_25 : std_logic;
	signal N8_1_26 : std_logic;
	signal N8_2_25 : std_logic;
	signal N8_3_26 : std_logic;
	signal N8_0_26 : std_logic;
	signal N8_1_27 : std_logic;
	signal N8_2_26 : std_logic;
	signal N8_3_27 : std_logic;
	signal N8_0_27 : std_logic;
	signal N8_1_28 : std_logic;
	signal N8_2_27 : std_logic;
	signal N8_3_28 : std_logic;
	signal N8_0_28 : std_logic;
	signal N8_1_29 : std_logic;
	signal N8_2_28 : std_logic;
	signal N8_3_29 : std_logic;
	signal N8_0_29 : std_logic;
	signal N8_1_30 : std_logic;
	signal N8_2_29 : std_logic;
	signal N8_3_30 : std_logic;
	signal N8_0_30 : std_logic;
	signal N8_1_31 : std_logic;
	signal N8_2_30 : std_logic;
	signal N8_3_31 : std_logic;
	signal N8_0_31 : std_logic;
	signal N8_1_32 : std_logic;
	signal N8_2_31 : std_logic;
	signal N8_3_32 : std_logic;
	signal N8_0_32 : std_logic;
	signal N8_1_33 : std_logic;
	signal N8_2_32 : std_logic;
	signal N8_3_33 : std_logic;
	signal N8_0_33 : std_logic;
	signal N8_1_34 : std_logic;
	signal N8_2_33 : std_logic;
	signal N8_3_34 : std_logic;
	signal N8_0_34 : std_logic;
	signal N8_1_35 : std_logic;
	signal N8_2_34 : std_logic;
	signal N8_3_35 : std_logic;
	signal N8_0_35 : std_logic;
	signal N8_1_36 : std_logic;
	signal N8_2_35 : std_logic;
	signal N8_3_36 : std_logic;
	signal N8_0_36 : std_logic;
	signal N8_1_37 : std_logic;
	signal N8_2_36 : std_logic;
	signal N8_3_37 : std_logic;
	signal N8_0_37 : std_logic;
	signal N8_1_38 : std_logic;
	signal N8_2_37 : std_logic;
	signal N8_3_38 : std_logic;
	signal N8_0_38 : std_logic;
	signal N8_1_39 : std_logic;
	signal N8_2_38 : std_logic;
	signal N8_3_39 : std_logic;
	signal N8_0_39 : std_logic;
	signal N8_1_40 : std_logic;
	signal N8_2_39 : std_logic;
	signal N8_3_40 : std_logic;
	signal N8_0_40 : std_logic;
	signal N8_1_41 : std_logic;
	signal N8_2_40 : std_logic;
	signal N8_3_41 : std_logic;
	signal N8_0_41 : std_logic;
	signal N8_1_42 : std_logic;
	signal N8_2_41 : std_logic;
	signal N8_3_42 : std_logic;
	signal N8_0_42 : std_logic;
	signal N8_1_43 : std_logic;
	signal N8_2_42 : std_logic;
	signal N8_3_43 : std_logic;
	signal N8_0_43 : std_logic;
	signal N8_1_44 : std_logic;
	signal N8_2_43 : std_logic;
	signal N8_3_44 : std_logic;
	signal N8_0_44 : std_logic;
	signal N8_1_45 : std_logic;
	signal N8_2_44 : std_logic;
	signal N8_3_45 : std_logic;
	signal N8_0_45 : std_logic;
	signal N8_1_46 : std_logic;
	signal N8_2_45 : std_logic;
	signal N8_3_46 : std_logic;
	signal N8_0_46 : std_logic;
	signal N8_1_47 : std_logic;
	signal N8_2_46 : std_logic;
	signal N8_3_47 : std_logic;
	signal N8_0_47 : std_logic;
	signal N8_1_48 : std_logic;
	signal N8_2_47 : std_logic;
	signal N8_3_48 : std_logic;
	signal N8_0_48 : std_logic;
	signal N8_1_49 : std_logic;
	signal N8_2_48 : std_logic;
	signal N8_3_49 : std_logic;
	signal N8_0_49 : std_logic;
	signal N8_1_50 : std_logic;
	signal N8_2_49 : std_logic;
	signal N8_3_50 : std_logic;
	signal N8_0_50 : std_logic;
	signal N8_1_51 : std_logic;
	signal N8_2_50 : std_logic;
	signal N8_3_51 : std_logic;
	signal N8_0_51 : std_logic;
	signal N8_1_52 : std_logic;
	signal N8_2_51 : std_logic;
	signal N8_3_52 : std_logic;
	signal N8_0_52 : std_logic;
	signal N8_1_53 : std_logic;
	signal N8_2_52 : std_logic;
	signal N8_3_53 : std_logic;
	signal N8_0_53 : std_logic;
	signal N8_1_54 : std_logic;
	signal N8_2_53 : std_logic;
	signal N8_3_54 : std_logic;
	signal N8_0_54 : std_logic;
	signal N8_1_55 : std_logic;
	signal N8_2_54 : std_logic;
	signal N8_3_55 : std_logic;
	signal N8_0_55 : std_logic;
	signal N8_1_56 : std_logic;
	signal N8_2_55 : std_logic;
	signal N8_3_56 : std_logic;
	signal N8_0_56 : std_logic;
	signal N8_1_57 : std_logic;
	signal N8_2_56 : std_logic;
	signal N8_3_57 : std_logic;
	signal N8_0_57 : std_logic;
	signal N8_1_58 : std_logic;
	signal N8_2_57 : std_logic;
	signal N8_3_58 : std_logic;
	signal N8_0_58 : std_logic;
	signal N8_1_59 : std_logic;
	signal N8_2_58 : std_logic;
	signal N8_3_59 : std_logic;
	signal N8_0_59 : std_logic;
	signal N8_1_60 : std_logic;
	signal N8_2_59 : std_logic;
	signal N8_3_60 : std_logic;
	signal N8_0_60 : std_logic;
	signal N8_1_61 : std_logic;
	signal N8_2_60 : std_logic;
	signal N8_3_61 : std_logic;
	signal N8_0_61 : std_logic;
	signal N8_1_62 : std_logic;
	signal N8_2_61 : std_logic;
	signal N8_3_62 : std_logic;
	signal N8_0_62 : std_logic;
	signal N8_1_63 : std_logic;
	signal N8_2_62 : std_logic;
	signal N8_3_63 : std_logic;
	signal N8_0_63 : std_logic;
	signal N8_1_64 : std_logic;
	signal N8_2_63 : std_logic;
	signal N8_3_64 : std_logic;
	signal N8_0_64 : std_logic;
	signal N8_1_65 : std_logic;
	signal N8_2_64 : std_logic;
	signal N8_3_65 : std_logic;
	signal N8_0_65 : std_logic;
	signal N8_1_66 : std_logic;
	signal N8_2_65 : std_logic;
	signal N8_3_66 : std_logic;
	signal N8_0_66 : std_logic;
	signal N8_1_67 : std_logic;
	signal N8_2_66 : std_logic;
	signal N8_3_67 : std_logic;
	signal N8_0_67 : std_logic;
	signal N8_1_68 : std_logic;
	signal N8_2_67 : std_logic;
	signal N8_3_68 : std_logic;
	signal N8_0_68 : std_logic;
	signal N8_1_69 : std_logic;
	signal N8_2_68 : std_logic;
	signal N8_3_69 : std_logic;
	signal N8_0_69 : std_logic;
	signal N8_1_70 : std_logic;
	signal N8_2_69 : std_logic;
	signal N8_3_70 : std_logic;
	signal N8_0_70 : std_logic;
	signal N8_1_71 : std_logic;
	signal N8_2_70 : std_logic;
	signal N8_3_71 : std_logic;
	signal N8_0_71 : std_logic;
	signal N8_1_72 : std_logic;
	signal N8_2_71 : std_logic;
	signal N8_3_72 : std_logic;
	signal N8_0_72 : std_logic;
	signal N8_1_73 : std_logic;
	signal N8_2_72 : std_logic;
	signal N8_3_73 : std_logic;
	signal N8_0_73 : std_logic;
	signal N8_1_74 : std_logic;
	signal N8_2_73 : std_logic;
	signal N8_3_74 : std_logic;
	signal N8_0_74 : std_logic;
	signal N8_1_75 : std_logic;
	signal N8_2_74 : std_logic;
	signal N8_3_75 : std_logic;
	signal N8_0_75 : std_logic;
	signal N8_1_76 : std_logic;
	signal N8_2_75 : std_logic;
	signal N8_3_76 : std_logic;
	signal N8_0_76 : std_logic;
	signal N8_1_77 : std_logic;
	signal N8_2_76 : std_logic;
	signal N8_3_77 : std_logic;
	signal N8_0_77 : std_logic;
	signal N8_1_78 : std_logic;
	signal N8_2_77 : std_logic;
	signal N8_3_78 : std_logic;
	signal N8_0_78 : std_logic;
	signal N8_1_79 : std_logic;
	signal N8_2_78 : std_logic;
	signal N8_3_79 : std_logic;
	signal N8_0_79 : std_logic;
	signal N8_1_80 : std_logic;
	signal N8_2_79 : std_logic;
	signal N8_3_80 : std_logic;
	signal N8_0_80 : std_logic;
	signal N8_1_81 : std_logic;
	signal N8_2_80 : std_logic;
	signal N8_3_81 : std_logic;
	signal N8_0_81 : std_logic;
	signal N8_1_82 : std_logic;
	signal N8_2_81 : std_logic;
	signal N8_3_82 : std_logic;
	signal N8_0_82 : std_logic;
	signal N8_1_83 : std_logic;
	signal N8_2_82 : std_logic;
	signal N8_3_83 : std_logic;
	signal N8_0_83 : std_logic;
	signal N8_1_84 : std_logic;
	signal N8_2_83 : std_logic;
	signal N8_3_84 : std_logic;
	signal N8_0_84 : std_logic;
	signal N8_1_85 : std_logic;
	signal N8_2_84 : std_logic;
	signal N8_3_85 : std_logic;
	signal N8_0_85 : std_logic;
	signal N8_1_86 : std_logic;
	signal N8_2_85 : std_logic;
	signal N8_3_86 : std_logic;
	signal N8_0_86 : std_logic;
	signal N8_1_87 : std_logic;
	signal N8_2_86 : std_logic;
	signal N8_3_87 : std_logic;
	signal N8_0_87 : std_logic;
	signal N8_1_88 : std_logic;
	signal N8_2_87 : std_logic;
	signal N8_3_88 : std_logic;
	signal N8_0_88 : std_logic;
	signal N8_1_89 : std_logic;
	signal N8_2_88 : std_logic;
	signal N8_3_89 : std_logic;
	signal N8_0_89 : std_logic;
	signal N8_1_90 : std_logic;
	signal N8_2_89 : std_logic;
	signal N8_3_90 : std_logic;
	signal N8_0_90 : std_logic;
	signal N8_1_91 : std_logic;
	signal N8_2_90 : std_logic;
	signal N8_3_91 : std_logic;
	signal N8_0_91 : std_logic;
	signal N8_1_92 : std_logic;
	signal N8_2_91 : std_logic;
	signal N8_3_92 : std_logic;
	signal N8_0_92 : std_logic;
	signal N8_1_93 : std_logic;
	signal N8_2_92 : std_logic;
	signal N8_3_93 : std_logic;
	signal N8_0_93 : std_logic;
	signal N8_1_94 : std_logic;
	signal N8_2_93 : std_logic;
	signal N8_3_94 : std_logic;
	signal N8_0_94 : std_logic;
	signal N8_1_95 : std_logic;
	signal N8_2_94 : std_logic;
	signal N8_3_95 : std_logic;
	signal N8_0_95 : std_logic;
	signal N8_1_96 : std_logic;
	signal N8_2_95 : std_logic;
	signal N8_3_96 : std_logic;
	signal N8_0_96 : std_logic;
	signal N8_1_97 : std_logic;
	signal N8_2_96 : std_logic;
	signal N8_3_97 : std_logic;
	signal N8_0_97 : std_logic;
	signal N8_1_98 : std_logic;
	signal N8_2_97 : std_logic;
	signal N8_3_98 : std_logic;
	signal N8_0_98 : std_logic;
	signal N8_1_99 : std_logic;
	signal N8_2_98 : std_logic;
	signal N8_3_99 : std_logic;
	signal N8_0_99 : std_logic;
	signal N8_1_100 : std_logic;
	signal N8_2_99 : std_logic;
	signal N8_3_100 : std_logic;
	signal N8_0_100 : std_logic;
	signal N8_1_101 : std_logic;
	signal N8_2_100 : std_logic;
	signal N8_3_101 : std_logic;
	signal N8_0_101 : std_logic;
	signal N8_1_102 : std_logic;
	signal N9_0_3 : std_logic;
	signal N9_1_4 : std_logic;
	signal N9_0_4 : std_logic;
	signal N9_1_5 : std_logic;
	signal N9_0_5 : std_logic;
	signal N9_1_6 : std_logic;
	signal N9_0_6 : std_logic;
	signal N9_1_7 : std_logic;
	signal N9_0_7 : std_logic;
	signal N9_1_8 : std_logic;
	signal N9_0_8 : std_logic;
	signal N9_1_9 : std_logic;
	signal N9_0_9 : std_logic;
	signal N9_1_10 : std_logic;
	signal N9_0_10 : std_logic;
	signal N9_1_11 : std_logic;
	signal N9_0_11 : std_logic;
	signal N9_1_12 : std_logic;
	signal N9_0_12 : std_logic;
	signal N9_1_13 : std_logic;
	signal N9_0_13 : std_logic;
	signal N9_1_14 : std_logic;
	signal N9_0_14 : std_logic;
	signal N9_1_15 : std_logic;
	signal N9_0_15 : std_logic;
	signal N9_1_16 : std_logic;
	signal N9_0_16 : std_logic;
	signal N9_1_17 : std_logic;
	signal N9_0_17 : std_logic;
	signal N9_1_18 : std_logic;
	signal N9_0_18 : std_logic;
	signal N9_1_19 : std_logic;
	signal N9_0_19 : std_logic;
	signal N9_1_20 : std_logic;
	signal N9_0_20 : std_logic;
	signal N9_1_21 : std_logic;
	signal N9_0_21 : std_logic;
	signal N9_1_22 : std_logic;
	signal N9_0_22 : std_logic;
	signal N9_1_23 : std_logic;
	signal N9_0_23 : std_logic;
	signal N9_1_24 : std_logic;
	signal N9_0_24 : std_logic;
	signal N9_1_25 : std_logic;
	signal N9_0_25 : std_logic;
	signal N9_1_26 : std_logic;
	signal N9_0_26 : std_logic;
	signal N9_1_27 : std_logic;
	signal N9_0_27 : std_logic;
	signal N9_1_28 : std_logic;
	signal N9_0_28 : std_logic;
	signal N9_1_29 : std_logic;
	signal N9_0_29 : std_logic;
	signal N9_1_30 : std_logic;
	signal N9_0_30 : std_logic;
	signal N9_1_31 : std_logic;
	signal N9_0_31 : std_logic;
	signal N9_1_32 : std_logic;
	signal N9_0_32 : std_logic;
	signal N9_1_33 : std_logic;
	signal N9_0_33 : std_logic;
	signal N9_1_34 : std_logic;
	signal N9_0_34 : std_logic;
	signal N9_1_35 : std_logic;
	signal N9_0_35 : std_logic;
	signal N9_1_36 : std_logic;
	signal N9_0_36 : std_logic;
	signal N9_1_37 : std_logic;
	signal N9_0_37 : std_logic;
	signal N9_1_38 : std_logic;
	signal N9_0_38 : std_logic;
	signal N9_1_39 : std_logic;
	signal N9_0_39 : std_logic;
	signal N9_1_40 : std_logic;
	signal N9_0_40 : std_logic;
	signal N9_1_41 : std_logic;
	signal N9_0_41 : std_logic;
	signal N9_1_42 : std_logic;
	signal N9_0_42 : std_logic;
	signal N9_1_43 : std_logic;
	signal N9_0_43 : std_logic;
	signal N9_1_44 : std_logic;
	signal N9_0_44 : std_logic;
	signal N9_1_45 : std_logic;
	signal N9_0_45 : std_logic;
	signal N9_1_46 : std_logic;
	signal N9_0_46 : std_logic;
	signal N9_1_47 : std_logic;
	signal N9_0_47 : std_logic;
	signal N9_1_48 : std_logic;
	signal N9_0_48 : std_logic;
	signal N9_1_49 : std_logic;
	signal N9_0_49 : std_logic;
	signal N9_1_50 : std_logic;
	signal N9_0_50 : std_logic;
	signal N9_1_51 : std_logic;
	signal N9_0_51 : std_logic;
	signal N9_1_52 : std_logic;
	signal N9_0_52 : std_logic;
	signal N9_1_53 : std_logic;
	signal N9_0_53 : std_logic;
	signal N9_1_54 : std_logic;
	signal N9_0_54 : std_logic;
	signal N9_1_55 : std_logic;
	signal N9_0_55 : std_logic;
	signal N9_1_56 : std_logic;
	signal N9_0_56 : std_logic;
	signal N9_1_57 : std_logic;
	signal N9_0_57 : std_logic;
	signal N9_1_58 : std_logic;
	signal N9_0_58 : std_logic;
	signal N9_1_59 : std_logic;
	signal N9_0_59 : std_logic;
	signal N9_1_60 : std_logic;
	signal N9_0_60 : std_logic;
	signal N9_1_61 : std_logic;
	signal N9_0_61 : std_logic;
	signal N9_1_62 : std_logic;
	signal N9_0_62 : std_logic;
	signal N9_1_63 : std_logic;
	signal N9_0_63 : std_logic;
	signal N9_1_64 : std_logic;
	signal N9_0_64 : std_logic;
	signal N9_1_65 : std_logic;
	signal N9_0_65 : std_logic;
	signal N9_1_66 : std_logic;
	signal N9_0_66 : std_logic;
	signal N9_1_67 : std_logic;
	signal N9_0_67 : std_logic;
	signal N9_1_68 : std_logic;
	signal N9_0_68 : std_logic;
	signal N9_1_69 : std_logic;
	signal N9_0_69 : std_logic;
	signal N9_1_70 : std_logic;
	signal N9_0_70 : std_logic;
	signal N9_1_71 : std_logic;
	signal N9_0_71 : std_logic;
	signal N9_1_72 : std_logic;
	signal N9_0_72 : std_logic;
	signal N9_1_73 : std_logic;
	signal N9_0_73 : std_logic;
	signal N9_1_74 : std_logic;
	signal N9_0_74 : std_logic;
	signal N9_1_75 : std_logic;
	signal N9_0_75 : std_logic;
	signal N9_1_76 : std_logic;
	signal N9_0_76 : std_logic;
	signal N9_1_77 : std_logic;
	signal N9_0_77 : std_logic;
	signal N9_1_78 : std_logic;
	signal N9_0_78 : std_logic;
	signal N9_1_79 : std_logic;
	signal N9_0_79 : std_logic;
	signal N9_1_80 : std_logic;
	signal N9_0_80 : std_logic;
	signal N9_1_81 : std_logic;
	signal N9_0_81 : std_logic;
	signal N9_1_82 : std_logic;
	signal N9_0_82 : std_logic;
	signal N9_1_83 : std_logic;
	signal N9_0_83 : std_logic;
	signal N9_1_84 : std_logic;
	signal N9_0_84 : std_logic;
	signal N9_1_85 : std_logic;
	signal N9_0_85 : std_logic;
	signal N9_1_86 : std_logic;
	signal N9_0_86 : std_logic;
	signal N9_1_87 : std_logic;
	signal N9_0_87 : std_logic;
	signal N9_1_88 : std_logic;
	signal N9_0_88 : std_logic;
	signal N9_1_89 : std_logic;
	signal N9_0_89 : std_logic;
	signal N9_1_90 : std_logic;
	signal N9_0_90 : std_logic;
	signal N9_1_91 : std_logic;
	signal N9_0_91 : std_logic;
	signal N9_1_92 : std_logic;
	signal N9_0_92 : std_logic;
	signal N9_1_93 : std_logic;
	signal N9_0_93 : std_logic;
	signal N9_1_94 : std_logic;
	signal N9_0_94 : std_logic;
	signal N9_1_95 : std_logic;
	signal N9_0_95 : std_logic;
	signal N9_1_96 : std_logic;
	signal N9_0_96 : std_logic;
	signal N9_1_97 : std_logic;
	signal N9_0_97 : std_logic;
	signal N9_1_98 : std_logic;
	signal N9_0_98 : std_logic;
	signal N9_1_99 : std_logic;
	signal N9_0_99 : std_logic;
	signal N9_1_100 : std_logic;
	signal N9_0_100 : std_logic;
	signal N9_1_101 : std_logic;
	signal N9_0_101 : std_logic;
	signal N9_1_102 : std_logic;
	signal N9_0_102 : std_logic;
	signal N9_1_103 : std_logic;
	signal N10_0_2 : std_logic;
	signal N10_1_3 : std_logic;
	signal N10_0_3 : std_logic;
	signal N10_1_4 : std_logic;
	signal N10_0_4 : std_logic;
	signal N10_1_5 : std_logic;
	signal N10_0_5 : std_logic;
	signal N10_1_6 : std_logic;
	signal N10_0_6 : std_logic;
	signal N10_1_7 : std_logic;
	signal N10_0_7 : std_logic;
	signal N10_1_8 : std_logic;
	signal N10_0_8 : std_logic;
	signal N10_1_9 : std_logic;
	signal N10_0_9 : std_logic;
	signal N10_1_10 : std_logic;
	signal N10_0_10 : std_logic;
	signal N10_1_11 : std_logic;
	signal N10_0_11 : std_logic;
	signal N10_1_12 : std_logic;
	signal N10_0_12 : std_logic;
	signal N10_1_13 : std_logic;
	signal N10_0_13 : std_logic;
	signal N10_1_14 : std_logic;
	signal N10_0_14 : std_logic;
	signal N10_1_15 : std_logic;
	signal N10_0_15 : std_logic;
	signal N10_1_16 : std_logic;
	signal N10_0_16 : std_logic;
	signal N10_1_17 : std_logic;
	signal N10_0_17 : std_logic;
	signal N10_1_18 : std_logic;
	signal N10_0_18 : std_logic;
	signal N10_1_19 : std_logic;
	signal N10_0_19 : std_logic;
	signal N10_1_20 : std_logic;
	signal N10_0_20 : std_logic;
	signal N10_1_21 : std_logic;
	signal N10_0_21 : std_logic;
	signal N10_1_22 : std_logic;
	signal N10_0_22 : std_logic;
	signal N10_1_23 : std_logic;
	signal N10_0_23 : std_logic;
	signal N10_1_24 : std_logic;
	signal N10_0_24 : std_logic;
	signal N10_1_25 : std_logic;
	signal N10_0_25 : std_logic;
	signal N10_1_26 : std_logic;
	signal N10_0_26 : std_logic;
	signal N10_1_27 : std_logic;
	signal N10_0_27 : std_logic;
	signal N10_1_28 : std_logic;
	signal N10_0_28 : std_logic;
	signal N10_1_29 : std_logic;
	signal N10_0_29 : std_logic;
	signal N10_1_30 : std_logic;
	signal N10_0_30 : std_logic;
	signal N10_1_31 : std_logic;
	signal N10_0_31 : std_logic;
	signal N10_1_32 : std_logic;
	signal N10_0_32 : std_logic;
	signal N10_1_33 : std_logic;
	signal N10_0_33 : std_logic;
	signal N10_1_34 : std_logic;
	signal N10_0_34 : std_logic;
	signal N10_1_35 : std_logic;
	signal N10_0_35 : std_logic;
	signal N10_1_36 : std_logic;
	signal N10_0_36 : std_logic;
	signal N10_1_37 : std_logic;
	signal N10_0_37 : std_logic;
	signal N10_1_38 : std_logic;
	signal N10_0_38 : std_logic;
	signal N10_1_39 : std_logic;
	signal N10_0_39 : std_logic;
	signal N10_1_40 : std_logic;
	signal N10_0_40 : std_logic;
	signal N10_1_41 : std_logic;
	signal N10_0_41 : std_logic;
	signal N10_1_42 : std_logic;
	signal N10_0_42 : std_logic;
	signal N10_1_43 : std_logic;
	signal N10_0_43 : std_logic;
	signal N10_1_44 : std_logic;
	signal N10_0_44 : std_logic;
	signal N10_1_45 : std_logic;
	signal N10_0_45 : std_logic;
	signal N10_1_46 : std_logic;
	signal N10_0_46 : std_logic;
	signal N10_1_47 : std_logic;
	signal N10_0_47 : std_logic;
	signal N10_1_48 : std_logic;
	signal N10_0_48 : std_logic;
	signal N10_1_49 : std_logic;
	signal N10_0_49 : std_logic;
	signal N10_1_50 : std_logic;
	signal N10_0_50 : std_logic;
	signal N10_1_51 : std_logic;
	signal N10_0_51 : std_logic;
	signal N10_1_52 : std_logic;
	signal N10_0_52 : std_logic;
	signal N10_1_53 : std_logic;
	signal N10_0_53 : std_logic;
	signal N10_1_54 : std_logic;
	signal N10_0_54 : std_logic;
	signal N10_1_55 : std_logic;
	signal N10_0_55 : std_logic;
	signal N10_1_56 : std_logic;
	signal N10_0_56 : std_logic;
	signal N10_1_57 : std_logic;
	signal N10_0_57 : std_logic;
	signal N10_1_58 : std_logic;
	signal N10_0_58 : std_logic;
	signal N10_1_59 : std_logic;
	signal N10_0_59 : std_logic;
	signal N10_1_60 : std_logic;
	signal N10_0_60 : std_logic;
	signal N10_1_61 : std_logic;
	signal N10_0_61 : std_logic;
	signal N10_1_62 : std_logic;
	signal N10_0_62 : std_logic;
	signal N10_1_63 : std_logic;
	signal N10_0_63 : std_logic;
	signal N10_1_64 : std_logic;
	signal N10_0_64 : std_logic;
	signal N10_1_65 : std_logic;
	signal N10_0_65 : std_logic;
	signal N10_1_66 : std_logic;
	signal N10_0_66 : std_logic;
	signal N10_1_67 : std_logic;
	signal N10_0_67 : std_logic;
	signal N10_1_68 : std_logic;
	signal N10_0_68 : std_logic;
	signal N10_1_69 : std_logic;
	signal N10_0_69 : std_logic;
	signal N10_1_70 : std_logic;
	signal N10_0_70 : std_logic;
	signal N10_1_71 : std_logic;
	signal N10_0_71 : std_logic;
	signal N10_1_72 : std_logic;
	signal N10_0_72 : std_logic;
	signal N10_1_73 : std_logic;
	signal N10_0_73 : std_logic;
	signal N10_1_74 : std_logic;
	signal N10_0_74 : std_logic;
	signal N10_1_75 : std_logic;
	signal N10_0_75 : std_logic;
	signal N10_1_76 : std_logic;
	signal N10_0_76 : std_logic;
	signal N10_1_77 : std_logic;
	signal N10_0_77 : std_logic;
	signal N10_1_78 : std_logic;
	signal N10_0_78 : std_logic;
	signal N10_1_79 : std_logic;
	signal N10_0_79 : std_logic;
	signal N10_1_80 : std_logic;
	signal N10_0_80 : std_logic;
	signal N10_1_81 : std_logic;
	signal N10_0_81 : std_logic;
	signal N10_1_82 : std_logic;
	signal N10_0_82 : std_logic;
	signal N10_1_83 : std_logic;
	signal N10_0_83 : std_logic;
	signal N10_1_84 : std_logic;
	signal N10_0_84 : std_logic;
	signal N10_1_85 : std_logic;
	signal N10_0_85 : std_logic;
	signal N10_1_86 : std_logic;
	signal N10_0_86 : std_logic;
	signal N10_1_87 : std_logic;
	signal N10_0_87 : std_logic;
	signal N10_1_88 : std_logic;
	signal N10_0_88 : std_logic;
	signal N10_1_89 : std_logic;
	signal N10_0_89 : std_logic;
	signal N10_1_90 : std_logic;
	signal N10_0_90 : std_logic;
	signal N10_1_91 : std_logic;
	signal N10_0_91 : std_logic;
	signal N10_1_92 : std_logic;
	signal N10_0_92 : std_logic;
	signal N10_1_93 : std_logic;
	signal N10_0_93 : std_logic;
	signal N10_1_94 : std_logic;
	signal N10_0_94 : std_logic;
	signal N10_1_95 : std_logic;
	signal N10_0_95 : std_logic;
	signal N10_1_96 : std_logic;
	signal N10_0_96 : std_logic;
	signal N10_1_97 : std_logic;
	signal N10_0_97 : std_logic;
	signal N10_1_98 : std_logic;
	signal N10_0_98 : std_logic;
	signal N10_1_99 : std_logic;
	signal N10_0_99 : std_logic;
	signal N10_1_100 : std_logic;
	signal N10_0_100 : std_logic;
	signal N10_1_101 : std_logic;
	signal N10_0_101 : std_logic;
	signal N10_1_102 : std_logic;
	signal N10_0_102 : std_logic;
	signal N10_1_103 : std_logic;
	signal N10_0_103 : std_logic;
	signal N10_1_104 : std_logic;


begin
-- generate the partial products.
	-- signal N0_0_0 : std_logic;
	PP1 : and2 port map (X(0), Y(0), N0_0_0);
	-- signal N0_0_1 : std_logic;
	PP2 : and2 port map (X(1), Y(0), N0_0_1);
	-- signal N0_0_2 : std_logic;
	PP3 : and2 port map (X(2), Y(0), N0_0_2);
	-- signal N0_0_3 : std_logic;
	PP4 : and2 port map (X(3), Y(0), N0_0_3);
	-- signal N0_0_4 : std_logic;
	PP5 : and2 port map (X(4), Y(0), N0_0_4);
	-- signal N0_0_5 : std_logic;
	PP6 : and2 port map (X(5), Y(0), N0_0_5);
	-- signal N0_0_6 : std_logic;
	PP7 : and2 port map (X(6), Y(0), N0_0_6);
	-- signal N0_0_7 : std_logic;
	PP8 : and2 port map (X(7), Y(0), N0_0_7);
	-- signal N0_0_8 : std_logic;
	PP9 : and2 port map (X(8), Y(0), N0_0_8);
	-- signal N0_0_9 : std_logic;
	PP10 : and2 port map (X(9), Y(0), N0_0_9);
	-- signal N0_0_10 : std_logic;
	PP11 : and2 port map (X(10), Y(0), N0_0_10);
	-- signal N0_0_11 : std_logic;
	PP12 : and2 port map (X(11), Y(0), N0_0_11);
	-- signal N0_0_12 : std_logic;
	PP13 : and2 port map (X(12), Y(0), N0_0_12);
	-- signal N0_0_13 : std_logic;
	PP14 : and2 port map (X(13), Y(0), N0_0_13);
	-- signal N0_0_14 : std_logic;
	PP15 : and2 port map (X(14), Y(0), N0_0_14);
	-- signal N0_0_15 : std_logic;
	PP16 : and2 port map (X(15), Y(0), N0_0_15);
	-- signal N0_0_16 : std_logic;
	PP17 : and2 port map (X(16), Y(0), N0_0_16);
	-- signal N0_0_17 : std_logic;
	PP18 : and2 port map (X(17), Y(0), N0_0_17);
	-- signal N0_0_18 : std_logic;
	PP19 : and2 port map (X(18), Y(0), N0_0_18);
	-- signal N0_0_19 : std_logic;
	PP20 : and2 port map (X(19), Y(0), N0_0_19);
	-- signal N0_0_20 : std_logic;
	PP21 : and2 port map (X(20), Y(0), N0_0_20);
	-- signal N0_0_21 : std_logic;
	PP22 : and2 port map (X(21), Y(0), N0_0_21);
	-- signal N0_0_22 : std_logic;
	PP23 : and2 port map (X(22), Y(0), N0_0_22);
	-- signal N0_0_23 : std_logic;
	PP24 : and2 port map (X(23), Y(0), N0_0_23);
	-- signal N0_0_24 : std_logic;
	PP25 : and2 port map (X(24), Y(0), N0_0_24);
	-- signal N0_0_25 : std_logic;
	PP26 : and2 port map (X(25), Y(0), N0_0_25);
	-- signal N0_0_26 : std_logic;
	PP27 : and2 port map (X(26), Y(0), N0_0_26);
	-- signal N0_0_27 : std_logic;
	PP28 : and2 port map (X(27), Y(0), N0_0_27);
	-- signal N0_0_28 : std_logic;
	PP29 : and2 port map (X(28), Y(0), N0_0_28);
	-- signal N0_0_29 : std_logic;
	PP30 : and2 port map (X(29), Y(0), N0_0_29);
	-- signal N0_0_30 : std_logic;
	PP31 : and2 port map (X(30), Y(0), N0_0_30);
	-- signal N0_0_31 : std_logic;
	PP32 : and2 port map (X(31), Y(0), N0_0_31);
	-- signal N0_0_32 : std_logic;
	PP33 : and2 port map (X(32), Y(0), N0_0_32);
	-- signal N0_0_33 : std_logic;
	PP34 : and2 port map (X(33), Y(0), N0_0_33);
	-- signal N0_0_34 : std_logic;
	PP35 : and2 port map (X(34), Y(0), N0_0_34);
	-- signal N0_0_35 : std_logic;
	PP36 : and2 port map (X(35), Y(0), N0_0_35);
	-- signal N0_0_36 : std_logic;
	PP37 : and2 port map (X(36), Y(0), N0_0_36);
	-- signal N0_0_37 : std_logic;
	PP38 : and2 port map (X(37), Y(0), N0_0_37);
	-- signal N0_0_38 : std_logic;
	PP39 : and2 port map (X(38), Y(0), N0_0_38);
	-- signal N0_0_39 : std_logic;
	PP40 : and2 port map (X(39), Y(0), N0_0_39);
	-- signal N0_0_40 : std_logic;
	PP41 : and2 port map (X(40), Y(0), N0_0_40);
	-- signal N0_0_41 : std_logic;
	PP42 : and2 port map (X(41), Y(0), N0_0_41);
	-- signal N0_0_42 : std_logic;
	PP43 : and2 port map (X(42), Y(0), N0_0_42);
	-- signal N0_0_43 : std_logic;
	PP44 : and2 port map (X(43), Y(0), N0_0_43);
	-- signal N0_0_44 : std_logic;
	PP45 : and2 port map (X(44), Y(0), N0_0_44);
	-- signal N0_0_45 : std_logic;
	PP46 : and2 port map (X(45), Y(0), N0_0_45);
	-- signal N0_0_46 : std_logic;
	PP47 : and2 port map (X(46), Y(0), N0_0_46);
	-- signal N0_0_47 : std_logic;
	PP48 : and2 port map (X(47), Y(0), N0_0_47);
	-- signal N0_0_48 : std_logic;
	PP49 : and2 port map (X(48), Y(0), N0_0_48);
	-- signal N0_0_49 : std_logic;
	PP50 : and2 port map (X(49), Y(0), N0_0_49);
	-- signal N0_0_50 : std_logic;
	PP51 : and2 port map (X(50), Y(0), N0_0_50);
	-- signal N0_0_51 : std_logic;
	PP52 : and2 port map (X(51), Y(0), N0_0_51);
	-- signal N0_0_52 : std_logic;
	PP53 : and2 port map ('1', Y(0), N0_0_52);
	-- signal N0_1_1 : std_logic;
	PP54 : and2 port map (X(0), Y(1), N0_1_1);
	-- signal N0_1_2 : std_logic;
	PP55 : and2 port map (X(1), Y(1), N0_1_2);
	-- signal N0_1_3 : std_logic;
	PP56 : and2 port map (X(2), Y(1), N0_1_3);
	-- signal N0_1_4 : std_logic;
	PP57 : and2 port map (X(3), Y(1), N0_1_4);
	-- signal N0_1_5 : std_logic;
	PP58 : and2 port map (X(4), Y(1), N0_1_5);
	-- signal N0_1_6 : std_logic;
	PP59 : and2 port map (X(5), Y(1), N0_1_6);
	-- signal N0_1_7 : std_logic;
	PP60 : and2 port map (X(6), Y(1), N0_1_7);
	-- signal N0_1_8 : std_logic;
	PP61 : and2 port map (X(7), Y(1), N0_1_8);
	-- signal N0_1_9 : std_logic;
	PP62 : and2 port map (X(8), Y(1), N0_1_9);
	-- signal N0_1_10 : std_logic;
	PP63 : and2 port map (X(9), Y(1), N0_1_10);
	-- signal N0_1_11 : std_logic;
	PP64 : and2 port map (X(10), Y(1), N0_1_11);
	-- signal N0_1_12 : std_logic;
	PP65 : and2 port map (X(11), Y(1), N0_1_12);
	-- signal N0_1_13 : std_logic;
	PP66 : and2 port map (X(12), Y(1), N0_1_13);
	-- signal N0_1_14 : std_logic;
	PP67 : and2 port map (X(13), Y(1), N0_1_14);
	-- signal N0_1_15 : std_logic;
	PP68 : and2 port map (X(14), Y(1), N0_1_15);
	-- signal N0_1_16 : std_logic;
	PP69 : and2 port map (X(15), Y(1), N0_1_16);
	-- signal N0_1_17 : std_logic;
	PP70 : and2 port map (X(16), Y(1), N0_1_17);
	-- signal N0_1_18 : std_logic;
	PP71 : and2 port map (X(17), Y(1), N0_1_18);
	-- signal N0_1_19 : std_logic;
	PP72 : and2 port map (X(18), Y(1), N0_1_19);
	-- signal N0_1_20 : std_logic;
	PP73 : and2 port map (X(19), Y(1), N0_1_20);
	-- signal N0_1_21 : std_logic;
	PP74 : and2 port map (X(20), Y(1), N0_1_21);
	-- signal N0_1_22 : std_logic;
	PP75 : and2 port map (X(21), Y(1), N0_1_22);
	-- signal N0_1_23 : std_logic;
	PP76 : and2 port map (X(22), Y(1), N0_1_23);
	-- signal N0_1_24 : std_logic;
	PP77 : and2 port map (X(23), Y(1), N0_1_24);
	-- signal N0_1_25 : std_logic;
	PP78 : and2 port map (X(24), Y(1), N0_1_25);
	-- signal N0_1_26 : std_logic;
	PP79 : and2 port map (X(25), Y(1), N0_1_26);
	-- signal N0_1_27 : std_logic;
	PP80 : and2 port map (X(26), Y(1), N0_1_27);
	-- signal N0_1_28 : std_logic;
	PP81 : and2 port map (X(27), Y(1), N0_1_28);
	-- signal N0_1_29 : std_logic;
	PP82 : and2 port map (X(28), Y(1), N0_1_29);
	-- signal N0_1_30 : std_logic;
	PP83 : and2 port map (X(29), Y(1), N0_1_30);
	-- signal N0_1_31 : std_logic;
	PP84 : and2 port map (X(30), Y(1), N0_1_31);
	-- signal N0_1_32 : std_logic;
	PP85 : and2 port map (X(31), Y(1), N0_1_32);
	-- signal N0_1_33 : std_logic;
	PP86 : and2 port map (X(32), Y(1), N0_1_33);
	-- signal N0_1_34 : std_logic;
	PP87 : and2 port map (X(33), Y(1), N0_1_34);
	-- signal N0_1_35 : std_logic;
	PP88 : and2 port map (X(34), Y(1), N0_1_35);
	-- signal N0_1_36 : std_logic;
	PP89 : and2 port map (X(35), Y(1), N0_1_36);
	-- signal N0_1_37 : std_logic;
	PP90 : and2 port map (X(36), Y(1), N0_1_37);
	-- signal N0_1_38 : std_logic;
	PP91 : and2 port map (X(37), Y(1), N0_1_38);
	-- signal N0_1_39 : std_logic;
	PP92 : and2 port map (X(38), Y(1), N0_1_39);
	-- signal N0_1_40 : std_logic;
	PP93 : and2 port map (X(39), Y(1), N0_1_40);
	-- signal N0_1_41 : std_logic;
	PP94 : and2 port map (X(40), Y(1), N0_1_41);
	-- signal N0_1_42 : std_logic;
	PP95 : and2 port map (X(41), Y(1), N0_1_42);
	-- signal N0_1_43 : std_logic;
	PP96 : and2 port map (X(42), Y(1), N0_1_43);
	-- signal N0_1_44 : std_logic;
	PP97 : and2 port map (X(43), Y(1), N0_1_44);
	-- signal N0_1_45 : std_logic;
	PP98 : and2 port map (X(44), Y(1), N0_1_45);
	-- signal N0_1_46 : std_logic;
	PP99 : and2 port map (X(45), Y(1), N0_1_46);
	-- signal N0_1_47 : std_logic;
	PP100 : and2 port map (X(46), Y(1), N0_1_47);
	-- signal N0_1_48 : std_logic;
	PP101 : and2 port map (X(47), Y(1), N0_1_48);
	-- signal N0_1_49 : std_logic;
	PP102 : and2 port map (X(48), Y(1), N0_1_49);
	-- signal N0_1_50 : std_logic;
	PP103 : and2 port map (X(49), Y(1), N0_1_50);
	-- signal N0_1_51 : std_logic;
	PP104 : and2 port map (X(50), Y(1), N0_1_51);
	-- signal N0_1_52 : std_logic;
	PP105 : and2 port map (X(51), Y(1), N0_1_52);
	-- signal N0_1_53 : std_logic;
	PP106 : and2 port map ('1', Y(1), N0_1_53);
	-- signal N0_2_2 : std_logic;
	PP107 : and2 port map (X(0), Y(2), N0_2_2);
	-- signal N0_2_3 : std_logic;
	PP108 : and2 port map (X(1), Y(2), N0_2_3);
	-- signal N0_2_4 : std_logic;
	PP109 : and2 port map (X(2), Y(2), N0_2_4);
	-- signal N0_2_5 : std_logic;
	PP110 : and2 port map (X(3), Y(2), N0_2_5);
	-- signal N0_2_6 : std_logic;
	PP111 : and2 port map (X(4), Y(2), N0_2_6);
	-- signal N0_2_7 : std_logic;
	PP112 : and2 port map (X(5), Y(2), N0_2_7);
	-- signal N0_2_8 : std_logic;
	PP113 : and2 port map (X(6), Y(2), N0_2_8);
	-- signal N0_2_9 : std_logic;
	PP114 : and2 port map (X(7), Y(2), N0_2_9);
	-- signal N0_2_10 : std_logic;
	PP115 : and2 port map (X(8), Y(2), N0_2_10);
	-- signal N0_2_11 : std_logic;
	PP116 : and2 port map (X(9), Y(2), N0_2_11);
	-- signal N0_2_12 : std_logic;
	PP117 : and2 port map (X(10), Y(2), N0_2_12);
	-- signal N0_2_13 : std_logic;
	PP118 : and2 port map (X(11), Y(2), N0_2_13);
	-- signal N0_2_14 : std_logic;
	PP119 : and2 port map (X(12), Y(2), N0_2_14);
	-- signal N0_2_15 : std_logic;
	PP120 : and2 port map (X(13), Y(2), N0_2_15);
	-- signal N0_2_16 : std_logic;
	PP121 : and2 port map (X(14), Y(2), N0_2_16);
	-- signal N0_2_17 : std_logic;
	PP122 : and2 port map (X(15), Y(2), N0_2_17);
	-- signal N0_2_18 : std_logic;
	PP123 : and2 port map (X(16), Y(2), N0_2_18);
	-- signal N0_2_19 : std_logic;
	PP124 : and2 port map (X(17), Y(2), N0_2_19);
	-- signal N0_2_20 : std_logic;
	PP125 : and2 port map (X(18), Y(2), N0_2_20);
	-- signal N0_2_21 : std_logic;
	PP126 : and2 port map (X(19), Y(2), N0_2_21);
	-- signal N0_2_22 : std_logic;
	PP127 : and2 port map (X(20), Y(2), N0_2_22);
	-- signal N0_2_23 : std_logic;
	PP128 : and2 port map (X(21), Y(2), N0_2_23);
	-- signal N0_2_24 : std_logic;
	PP129 : and2 port map (X(22), Y(2), N0_2_24);
	-- signal N0_2_25 : std_logic;
	PP130 : and2 port map (X(23), Y(2), N0_2_25);
	-- signal N0_2_26 : std_logic;
	PP131 : and2 port map (X(24), Y(2), N0_2_26);
	-- signal N0_2_27 : std_logic;
	PP132 : and2 port map (X(25), Y(2), N0_2_27);
	-- signal N0_2_28 : std_logic;
	PP133 : and2 port map (X(26), Y(2), N0_2_28);
	-- signal N0_2_29 : std_logic;
	PP134 : and2 port map (X(27), Y(2), N0_2_29);
	-- signal N0_2_30 : std_logic;
	PP135 : and2 port map (X(28), Y(2), N0_2_30);
	-- signal N0_2_31 : std_logic;
	PP136 : and2 port map (X(29), Y(2), N0_2_31);
	-- signal N0_2_32 : std_logic;
	PP137 : and2 port map (X(30), Y(2), N0_2_32);
	-- signal N0_2_33 : std_logic;
	PP138 : and2 port map (X(31), Y(2), N0_2_33);
	-- signal N0_2_34 : std_logic;
	PP139 : and2 port map (X(32), Y(2), N0_2_34);
	-- signal N0_2_35 : std_logic;
	PP140 : and2 port map (X(33), Y(2), N0_2_35);
	-- signal N0_2_36 : std_logic;
	PP141 : and2 port map (X(34), Y(2), N0_2_36);
	-- signal N0_2_37 : std_logic;
	PP142 : and2 port map (X(35), Y(2), N0_2_37);
	-- signal N0_2_38 : std_logic;
	PP143 : and2 port map (X(36), Y(2), N0_2_38);
	-- signal N0_2_39 : std_logic;
	PP144 : and2 port map (X(37), Y(2), N0_2_39);
	-- signal N0_2_40 : std_logic;
	PP145 : and2 port map (X(38), Y(2), N0_2_40);
	-- signal N0_2_41 : std_logic;
	PP146 : and2 port map (X(39), Y(2), N0_2_41);
	-- signal N0_2_42 : std_logic;
	PP147 : and2 port map (X(40), Y(2), N0_2_42);
	-- signal N0_2_43 : std_logic;
	PP148 : and2 port map (X(41), Y(2), N0_2_43);
	-- signal N0_2_44 : std_logic;
	PP149 : and2 port map (X(42), Y(2), N0_2_44);
	-- signal N0_2_45 : std_logic;
	PP150 : and2 port map (X(43), Y(2), N0_2_45);
	-- signal N0_2_46 : std_logic;
	PP151 : and2 port map (X(44), Y(2), N0_2_46);
	-- signal N0_2_47 : std_logic;
	PP152 : and2 port map (X(45), Y(2), N0_2_47);
	-- signal N0_2_48 : std_logic;
	PP153 : and2 port map (X(46), Y(2), N0_2_48);
	-- signal N0_2_49 : std_logic;
	PP154 : and2 port map (X(47), Y(2), N0_2_49);
	-- signal N0_2_50 : std_logic;
	PP155 : and2 port map (X(48), Y(2), N0_2_50);
	-- signal N0_2_51 : std_logic;
	PP156 : and2 port map (X(49), Y(2), N0_2_51);
	-- signal N0_2_52 : std_logic;
	PP157 : and2 port map (X(50), Y(2), N0_2_52);
	-- signal N0_2_53 : std_logic;
	PP158 : and2 port map (X(51), Y(2), N0_2_53);
	-- signal N0_2_54 : std_logic;
	PP159 : and2 port map ('1', Y(2), N0_2_54);
	-- signal N0_3_3 : std_logic;
	PP160 : and2 port map (X(0), Y(3), N0_3_3);
	-- signal N0_3_4 : std_logic;
	PP161 : and2 port map (X(1), Y(3), N0_3_4);
	-- signal N0_3_5 : std_logic;
	PP162 : and2 port map (X(2), Y(3), N0_3_5);
	-- signal N0_3_6 : std_logic;
	PP163 : and2 port map (X(3), Y(3), N0_3_6);
	-- signal N0_3_7 : std_logic;
	PP164 : and2 port map (X(4), Y(3), N0_3_7);
	-- signal N0_3_8 : std_logic;
	PP165 : and2 port map (X(5), Y(3), N0_3_8);
	-- signal N0_3_9 : std_logic;
	PP166 : and2 port map (X(6), Y(3), N0_3_9);
	-- signal N0_3_10 : std_logic;
	PP167 : and2 port map (X(7), Y(3), N0_3_10);
	-- signal N0_3_11 : std_logic;
	PP168 : and2 port map (X(8), Y(3), N0_3_11);
	-- signal N0_3_12 : std_logic;
	PP169 : and2 port map (X(9), Y(3), N0_3_12);
	-- signal N0_3_13 : std_logic;
	PP170 : and2 port map (X(10), Y(3), N0_3_13);
	-- signal N0_3_14 : std_logic;
	PP171 : and2 port map (X(11), Y(3), N0_3_14);
	-- signal N0_3_15 : std_logic;
	PP172 : and2 port map (X(12), Y(3), N0_3_15);
	-- signal N0_3_16 : std_logic;
	PP173 : and2 port map (X(13), Y(3), N0_3_16);
	-- signal N0_3_17 : std_logic;
	PP174 : and2 port map (X(14), Y(3), N0_3_17);
	-- signal N0_3_18 : std_logic;
	PP175 : and2 port map (X(15), Y(3), N0_3_18);
	-- signal N0_3_19 : std_logic;
	PP176 : and2 port map (X(16), Y(3), N0_3_19);
	-- signal N0_3_20 : std_logic;
	PP177 : and2 port map (X(17), Y(3), N0_3_20);
	-- signal N0_3_21 : std_logic;
	PP178 : and2 port map (X(18), Y(3), N0_3_21);
	-- signal N0_3_22 : std_logic;
	PP179 : and2 port map (X(19), Y(3), N0_3_22);
	-- signal N0_3_23 : std_logic;
	PP180 : and2 port map (X(20), Y(3), N0_3_23);
	-- signal N0_3_24 : std_logic;
	PP181 : and2 port map (X(21), Y(3), N0_3_24);
	-- signal N0_3_25 : std_logic;
	PP182 : and2 port map (X(22), Y(3), N0_3_25);
	-- signal N0_3_26 : std_logic;
	PP183 : and2 port map (X(23), Y(3), N0_3_26);
	-- signal N0_3_27 : std_logic;
	PP184 : and2 port map (X(24), Y(3), N0_3_27);
	-- signal N0_3_28 : std_logic;
	PP185 : and2 port map (X(25), Y(3), N0_3_28);
	-- signal N0_3_29 : std_logic;
	PP186 : and2 port map (X(26), Y(3), N0_3_29);
	-- signal N0_3_30 : std_logic;
	PP187 : and2 port map (X(27), Y(3), N0_3_30);
	-- signal N0_3_31 : std_logic;
	PP188 : and2 port map (X(28), Y(3), N0_3_31);
	-- signal N0_3_32 : std_logic;
	PP189 : and2 port map (X(29), Y(3), N0_3_32);
	-- signal N0_3_33 : std_logic;
	PP190 : and2 port map (X(30), Y(3), N0_3_33);
	-- signal N0_3_34 : std_logic;
	PP191 : and2 port map (X(31), Y(3), N0_3_34);
	-- signal N0_3_35 : std_logic;
	PP192 : and2 port map (X(32), Y(3), N0_3_35);
	-- signal N0_3_36 : std_logic;
	PP193 : and2 port map (X(33), Y(3), N0_3_36);
	-- signal N0_3_37 : std_logic;
	PP194 : and2 port map (X(34), Y(3), N0_3_37);
	-- signal N0_3_38 : std_logic;
	PP195 : and2 port map (X(35), Y(3), N0_3_38);
	-- signal N0_3_39 : std_logic;
	PP196 : and2 port map (X(36), Y(3), N0_3_39);
	-- signal N0_3_40 : std_logic;
	PP197 : and2 port map (X(37), Y(3), N0_3_40);
	-- signal N0_3_41 : std_logic;
	PP198 : and2 port map (X(38), Y(3), N0_3_41);
	-- signal N0_3_42 : std_logic;
	PP199 : and2 port map (X(39), Y(3), N0_3_42);
	-- signal N0_3_43 : std_logic;
	PP200 : and2 port map (X(40), Y(3), N0_3_43);
	-- signal N0_3_44 : std_logic;
	PP201 : and2 port map (X(41), Y(3), N0_3_44);
	-- signal N0_3_45 : std_logic;
	PP202 : and2 port map (X(42), Y(3), N0_3_45);
	-- signal N0_3_46 : std_logic;
	PP203 : and2 port map (X(43), Y(3), N0_3_46);
	-- signal N0_3_47 : std_logic;
	PP204 : and2 port map (X(44), Y(3), N0_3_47);
	-- signal N0_3_48 : std_logic;
	PP205 : and2 port map (X(45), Y(3), N0_3_48);
	-- signal N0_3_49 : std_logic;
	PP206 : and2 port map (X(46), Y(3), N0_3_49);
	-- signal N0_3_50 : std_logic;
	PP207 : and2 port map (X(47), Y(3), N0_3_50);
	-- signal N0_3_51 : std_logic;
	PP208 : and2 port map (X(48), Y(3), N0_3_51);
	-- signal N0_3_52 : std_logic;
	PP209 : and2 port map (X(49), Y(3), N0_3_52);
	-- signal N0_3_53 : std_logic;
	PP210 : and2 port map (X(50), Y(3), N0_3_53);
	-- signal N0_3_54 : std_logic;
	PP211 : and2 port map (X(51), Y(3), N0_3_54);
	-- signal N0_3_55 : std_logic;
	PP212 : and2 port map ('1', Y(3), N0_3_55);
	-- signal N0_4_4 : std_logic;
	PP213 : and2 port map (X(0), Y(4), N0_4_4);
	-- signal N0_4_5 : std_logic;
	PP214 : and2 port map (X(1), Y(4), N0_4_5);
	-- signal N0_4_6 : std_logic;
	PP215 : and2 port map (X(2), Y(4), N0_4_6);
	-- signal N0_4_7 : std_logic;
	PP216 : and2 port map (X(3), Y(4), N0_4_7);
	-- signal N0_4_8 : std_logic;
	PP217 : and2 port map (X(4), Y(4), N0_4_8);
	-- signal N0_4_9 : std_logic;
	PP218 : and2 port map (X(5), Y(4), N0_4_9);
	-- signal N0_4_10 : std_logic;
	PP219 : and2 port map (X(6), Y(4), N0_4_10);
	-- signal N0_4_11 : std_logic;
	PP220 : and2 port map (X(7), Y(4), N0_4_11);
	-- signal N0_4_12 : std_logic;
	PP221 : and2 port map (X(8), Y(4), N0_4_12);
	-- signal N0_4_13 : std_logic;
	PP222 : and2 port map (X(9), Y(4), N0_4_13);
	-- signal N0_4_14 : std_logic;
	PP223 : and2 port map (X(10), Y(4), N0_4_14);
	-- signal N0_4_15 : std_logic;
	PP224 : and2 port map (X(11), Y(4), N0_4_15);
	-- signal N0_4_16 : std_logic;
	PP225 : and2 port map (X(12), Y(4), N0_4_16);
	-- signal N0_4_17 : std_logic;
	PP226 : and2 port map (X(13), Y(4), N0_4_17);
	-- signal N0_4_18 : std_logic;
	PP227 : and2 port map (X(14), Y(4), N0_4_18);
	-- signal N0_4_19 : std_logic;
	PP228 : and2 port map (X(15), Y(4), N0_4_19);
	-- signal N0_4_20 : std_logic;
	PP229 : and2 port map (X(16), Y(4), N0_4_20);
	-- signal N0_4_21 : std_logic;
	PP230 : and2 port map (X(17), Y(4), N0_4_21);
	-- signal N0_4_22 : std_logic;
	PP231 : and2 port map (X(18), Y(4), N0_4_22);
	-- signal N0_4_23 : std_logic;
	PP232 : and2 port map (X(19), Y(4), N0_4_23);
	-- signal N0_4_24 : std_logic;
	PP233 : and2 port map (X(20), Y(4), N0_4_24);
	-- signal N0_4_25 : std_logic;
	PP234 : and2 port map (X(21), Y(4), N0_4_25);
	-- signal N0_4_26 : std_logic;
	PP235 : and2 port map (X(22), Y(4), N0_4_26);
	-- signal N0_4_27 : std_logic;
	PP236 : and2 port map (X(23), Y(4), N0_4_27);
	-- signal N0_4_28 : std_logic;
	PP237 : and2 port map (X(24), Y(4), N0_4_28);
	-- signal N0_4_29 : std_logic;
	PP238 : and2 port map (X(25), Y(4), N0_4_29);
	-- signal N0_4_30 : std_logic;
	PP239 : and2 port map (X(26), Y(4), N0_4_30);
	-- signal N0_4_31 : std_logic;
	PP240 : and2 port map (X(27), Y(4), N0_4_31);
	-- signal N0_4_32 : std_logic;
	PP241 : and2 port map (X(28), Y(4), N0_4_32);
	-- signal N0_4_33 : std_logic;
	PP242 : and2 port map (X(29), Y(4), N0_4_33);
	-- signal N0_4_34 : std_logic;
	PP243 : and2 port map (X(30), Y(4), N0_4_34);
	-- signal N0_4_35 : std_logic;
	PP244 : and2 port map (X(31), Y(4), N0_4_35);
	-- signal N0_4_36 : std_logic;
	PP245 : and2 port map (X(32), Y(4), N0_4_36);
	-- signal N0_4_37 : std_logic;
	PP246 : and2 port map (X(33), Y(4), N0_4_37);
	-- signal N0_4_38 : std_logic;
	PP247 : and2 port map (X(34), Y(4), N0_4_38);
	-- signal N0_4_39 : std_logic;
	PP248 : and2 port map (X(35), Y(4), N0_4_39);
	-- signal N0_4_40 : std_logic;
	PP249 : and2 port map (X(36), Y(4), N0_4_40);
	-- signal N0_4_41 : std_logic;
	PP250 : and2 port map (X(37), Y(4), N0_4_41);
	-- signal N0_4_42 : std_logic;
	PP251 : and2 port map (X(38), Y(4), N0_4_42);
	-- signal N0_4_43 : std_logic;
	PP252 : and2 port map (X(39), Y(4), N0_4_43);
	-- signal N0_4_44 : std_logic;
	PP253 : and2 port map (X(40), Y(4), N0_4_44);
	-- signal N0_4_45 : std_logic;
	PP254 : and2 port map (X(41), Y(4), N0_4_45);
	-- signal N0_4_46 : std_logic;
	PP255 : and2 port map (X(42), Y(4), N0_4_46);
	-- signal N0_4_47 : std_logic;
	PP256 : and2 port map (X(43), Y(4), N0_4_47);
	-- signal N0_4_48 : std_logic;
	PP257 : and2 port map (X(44), Y(4), N0_4_48);
	-- signal N0_4_49 : std_logic;
	PP258 : and2 port map (X(45), Y(4), N0_4_49);
	-- signal N0_4_50 : std_logic;
	PP259 : and2 port map (X(46), Y(4), N0_4_50);
	-- signal N0_4_51 : std_logic;
	PP260 : and2 port map (X(47), Y(4), N0_4_51);
	-- signal N0_4_52 : std_logic;
	PP261 : and2 port map (X(48), Y(4), N0_4_52);
	-- signal N0_4_53 : std_logic;
	PP262 : and2 port map (X(49), Y(4), N0_4_53);
	-- signal N0_4_54 : std_logic;
	PP263 : and2 port map (X(50), Y(4), N0_4_54);
	-- signal N0_4_55 : std_logic;
	PP264 : and2 port map (X(51), Y(4), N0_4_55);
	-- signal N0_4_56 : std_logic;
	PP265 : and2 port map ('1', Y(4), N0_4_56);
	-- signal N0_5_5 : std_logic;
	PP266 : and2 port map (X(0), Y(5), N0_5_5);
	-- signal N0_5_6 : std_logic;
	PP267 : and2 port map (X(1), Y(5), N0_5_6);
	-- signal N0_5_7 : std_logic;
	PP268 : and2 port map (X(2), Y(5), N0_5_7);
	-- signal N0_5_8 : std_logic;
	PP269 : and2 port map (X(3), Y(5), N0_5_8);
	-- signal N0_5_9 : std_logic;
	PP270 : and2 port map (X(4), Y(5), N0_5_9);
	-- signal N0_5_10 : std_logic;
	PP271 : and2 port map (X(5), Y(5), N0_5_10);
	-- signal N0_5_11 : std_logic;
	PP272 : and2 port map (X(6), Y(5), N0_5_11);
	-- signal N0_5_12 : std_logic;
	PP273 : and2 port map (X(7), Y(5), N0_5_12);
	-- signal N0_5_13 : std_logic;
	PP274 : and2 port map (X(8), Y(5), N0_5_13);
	-- signal N0_5_14 : std_logic;
	PP275 : and2 port map (X(9), Y(5), N0_5_14);
	-- signal N0_5_15 : std_logic;
	PP276 : and2 port map (X(10), Y(5), N0_5_15);
	-- signal N0_5_16 : std_logic;
	PP277 : and2 port map (X(11), Y(5), N0_5_16);
	-- signal N0_5_17 : std_logic;
	PP278 : and2 port map (X(12), Y(5), N0_5_17);
	-- signal N0_5_18 : std_logic;
	PP279 : and2 port map (X(13), Y(5), N0_5_18);
	-- signal N0_5_19 : std_logic;
	PP280 : and2 port map (X(14), Y(5), N0_5_19);
	-- signal N0_5_20 : std_logic;
	PP281 : and2 port map (X(15), Y(5), N0_5_20);
	-- signal N0_5_21 : std_logic;
	PP282 : and2 port map (X(16), Y(5), N0_5_21);
	-- signal N0_5_22 : std_logic;
	PP283 : and2 port map (X(17), Y(5), N0_5_22);
	-- signal N0_5_23 : std_logic;
	PP284 : and2 port map (X(18), Y(5), N0_5_23);
	-- signal N0_5_24 : std_logic;
	PP285 : and2 port map (X(19), Y(5), N0_5_24);
	-- signal N0_5_25 : std_logic;
	PP286 : and2 port map (X(20), Y(5), N0_5_25);
	-- signal N0_5_26 : std_logic;
	PP287 : and2 port map (X(21), Y(5), N0_5_26);
	-- signal N0_5_27 : std_logic;
	PP288 : and2 port map (X(22), Y(5), N0_5_27);
	-- signal N0_5_28 : std_logic;
	PP289 : and2 port map (X(23), Y(5), N0_5_28);
	-- signal N0_5_29 : std_logic;
	PP290 : and2 port map (X(24), Y(5), N0_5_29);
	-- signal N0_5_30 : std_logic;
	PP291 : and2 port map (X(25), Y(5), N0_5_30);
	-- signal N0_5_31 : std_logic;
	PP292 : and2 port map (X(26), Y(5), N0_5_31);
	-- signal N0_5_32 : std_logic;
	PP293 : and2 port map (X(27), Y(5), N0_5_32);
	-- signal N0_5_33 : std_logic;
	PP294 : and2 port map (X(28), Y(5), N0_5_33);
	-- signal N0_5_34 : std_logic;
	PP295 : and2 port map (X(29), Y(5), N0_5_34);
	-- signal N0_5_35 : std_logic;
	PP296 : and2 port map (X(30), Y(5), N0_5_35);
	-- signal N0_5_36 : std_logic;
	PP297 : and2 port map (X(31), Y(5), N0_5_36);
	-- signal N0_5_37 : std_logic;
	PP298 : and2 port map (X(32), Y(5), N0_5_37);
	-- signal N0_5_38 : std_logic;
	PP299 : and2 port map (X(33), Y(5), N0_5_38);
	-- signal N0_5_39 : std_logic;
	PP300 : and2 port map (X(34), Y(5), N0_5_39);
	-- signal N0_5_40 : std_logic;
	PP301 : and2 port map (X(35), Y(5), N0_5_40);
	-- signal N0_5_41 : std_logic;
	PP302 : and2 port map (X(36), Y(5), N0_5_41);
	-- signal N0_5_42 : std_logic;
	PP303 : and2 port map (X(37), Y(5), N0_5_42);
	-- signal N0_5_43 : std_logic;
	PP304 : and2 port map (X(38), Y(5), N0_5_43);
	-- signal N0_5_44 : std_logic;
	PP305 : and2 port map (X(39), Y(5), N0_5_44);
	-- signal N0_5_45 : std_logic;
	PP306 : and2 port map (X(40), Y(5), N0_5_45);
	-- signal N0_5_46 : std_logic;
	PP307 : and2 port map (X(41), Y(5), N0_5_46);
	-- signal N0_5_47 : std_logic;
	PP308 : and2 port map (X(42), Y(5), N0_5_47);
	-- signal N0_5_48 : std_logic;
	PP309 : and2 port map (X(43), Y(5), N0_5_48);
	-- signal N0_5_49 : std_logic;
	PP310 : and2 port map (X(44), Y(5), N0_5_49);
	-- signal N0_5_50 : std_logic;
	PP311 : and2 port map (X(45), Y(5), N0_5_50);
	-- signal N0_5_51 : std_logic;
	PP312 : and2 port map (X(46), Y(5), N0_5_51);
	-- signal N0_5_52 : std_logic;
	PP313 : and2 port map (X(47), Y(5), N0_5_52);
	-- signal N0_5_53 : std_logic;
	PP314 : and2 port map (X(48), Y(5), N0_5_53);
	-- signal N0_5_54 : std_logic;
	PP315 : and2 port map (X(49), Y(5), N0_5_54);
	-- signal N0_5_55 : std_logic;
	PP316 : and2 port map (X(50), Y(5), N0_5_55);
	-- signal N0_5_56 : std_logic;
	PP317 : and2 port map (X(51), Y(5), N0_5_56);
	-- signal N0_5_57 : std_logic;
	PP318 : and2 port map ('1', Y(5), N0_5_57);
	-- signal N0_6_6 : std_logic;
	PP319 : and2 port map (X(0), Y(6), N0_6_6);
	-- signal N0_6_7 : std_logic;
	PP320 : and2 port map (X(1), Y(6), N0_6_7);
	-- signal N0_6_8 : std_logic;
	PP321 : and2 port map (X(2), Y(6), N0_6_8);
	-- signal N0_6_9 : std_logic;
	PP322 : and2 port map (X(3), Y(6), N0_6_9);
	-- signal N0_6_10 : std_logic;
	PP323 : and2 port map (X(4), Y(6), N0_6_10);
	-- signal N0_6_11 : std_logic;
	PP324 : and2 port map (X(5), Y(6), N0_6_11);
	-- signal N0_6_12 : std_logic;
	PP325 : and2 port map (X(6), Y(6), N0_6_12);
	-- signal N0_6_13 : std_logic;
	PP326 : and2 port map (X(7), Y(6), N0_6_13);
	-- signal N0_6_14 : std_logic;
	PP327 : and2 port map (X(8), Y(6), N0_6_14);
	-- signal N0_6_15 : std_logic;
	PP328 : and2 port map (X(9), Y(6), N0_6_15);
	-- signal N0_6_16 : std_logic;
	PP329 : and2 port map (X(10), Y(6), N0_6_16);
	-- signal N0_6_17 : std_logic;
	PP330 : and2 port map (X(11), Y(6), N0_6_17);
	-- signal N0_6_18 : std_logic;
	PP331 : and2 port map (X(12), Y(6), N0_6_18);
	-- signal N0_6_19 : std_logic;
	PP332 : and2 port map (X(13), Y(6), N0_6_19);
	-- signal N0_6_20 : std_logic;
	PP333 : and2 port map (X(14), Y(6), N0_6_20);
	-- signal N0_6_21 : std_logic;
	PP334 : and2 port map (X(15), Y(6), N0_6_21);
	-- signal N0_6_22 : std_logic;
	PP335 : and2 port map (X(16), Y(6), N0_6_22);
	-- signal N0_6_23 : std_logic;
	PP336 : and2 port map (X(17), Y(6), N0_6_23);
	-- signal N0_6_24 : std_logic;
	PP337 : and2 port map (X(18), Y(6), N0_6_24);
	-- signal N0_6_25 : std_logic;
	PP338 : and2 port map (X(19), Y(6), N0_6_25);
	-- signal N0_6_26 : std_logic;
	PP339 : and2 port map (X(20), Y(6), N0_6_26);
	-- signal N0_6_27 : std_logic;
	PP340 : and2 port map (X(21), Y(6), N0_6_27);
	-- signal N0_6_28 : std_logic;
	PP341 : and2 port map (X(22), Y(6), N0_6_28);
	-- signal N0_6_29 : std_logic;
	PP342 : and2 port map (X(23), Y(6), N0_6_29);
	-- signal N0_6_30 : std_logic;
	PP343 : and2 port map (X(24), Y(6), N0_6_30);
	-- signal N0_6_31 : std_logic;
	PP344 : and2 port map (X(25), Y(6), N0_6_31);
	-- signal N0_6_32 : std_logic;
	PP345 : and2 port map (X(26), Y(6), N0_6_32);
	-- signal N0_6_33 : std_logic;
	PP346 : and2 port map (X(27), Y(6), N0_6_33);
	-- signal N0_6_34 : std_logic;
	PP347 : and2 port map (X(28), Y(6), N0_6_34);
	-- signal N0_6_35 : std_logic;
	PP348 : and2 port map (X(29), Y(6), N0_6_35);
	-- signal N0_6_36 : std_logic;
	PP349 : and2 port map (X(30), Y(6), N0_6_36);
	-- signal N0_6_37 : std_logic;
	PP350 : and2 port map (X(31), Y(6), N0_6_37);
	-- signal N0_6_38 : std_logic;
	PP351 : and2 port map (X(32), Y(6), N0_6_38);
	-- signal N0_6_39 : std_logic;
	PP352 : and2 port map (X(33), Y(6), N0_6_39);
	-- signal N0_6_40 : std_logic;
	PP353 : and2 port map (X(34), Y(6), N0_6_40);
	-- signal N0_6_41 : std_logic;
	PP354 : and2 port map (X(35), Y(6), N0_6_41);
	-- signal N0_6_42 : std_logic;
	PP355 : and2 port map (X(36), Y(6), N0_6_42);
	-- signal N0_6_43 : std_logic;
	PP356 : and2 port map (X(37), Y(6), N0_6_43);
	-- signal N0_6_44 : std_logic;
	PP357 : and2 port map (X(38), Y(6), N0_6_44);
	-- signal N0_6_45 : std_logic;
	PP358 : and2 port map (X(39), Y(6), N0_6_45);
	-- signal N0_6_46 : std_logic;
	PP359 : and2 port map (X(40), Y(6), N0_6_46);
	-- signal N0_6_47 : std_logic;
	PP360 : and2 port map (X(41), Y(6), N0_6_47);
	-- signal N0_6_48 : std_logic;
	PP361 : and2 port map (X(42), Y(6), N0_6_48);
	-- signal N0_6_49 : std_logic;
	PP362 : and2 port map (X(43), Y(6), N0_6_49);
	-- signal N0_6_50 : std_logic;
	PP363 : and2 port map (X(44), Y(6), N0_6_50);
	-- signal N0_6_51 : std_logic;
	PP364 : and2 port map (X(45), Y(6), N0_6_51);
	-- signal N0_6_52 : std_logic;
	PP365 : and2 port map (X(46), Y(6), N0_6_52);
	-- signal N0_6_53 : std_logic;
	PP366 : and2 port map (X(47), Y(6), N0_6_53);
	-- signal N0_6_54 : std_logic;
	PP367 : and2 port map (X(48), Y(6), N0_6_54);
	-- signal N0_6_55 : std_logic;
	PP368 : and2 port map (X(49), Y(6), N0_6_55);
	-- signal N0_6_56 : std_logic;
	PP369 : and2 port map (X(50), Y(6), N0_6_56);
	-- signal N0_6_57 : std_logic;
	PP370 : and2 port map (X(51), Y(6), N0_6_57);
	-- signal N0_6_58 : std_logic;
	PP371 : and2 port map ('1', Y(6), N0_6_58);
	-- signal N0_7_7 : std_logic;
	PP372 : and2 port map (X(0), Y(7), N0_7_7);
	-- signal N0_7_8 : std_logic;
	PP373 : and2 port map (X(1), Y(7), N0_7_8);
	-- signal N0_7_9 : std_logic;
	PP374 : and2 port map (X(2), Y(7), N0_7_9);
	-- signal N0_7_10 : std_logic;
	PP375 : and2 port map (X(3), Y(7), N0_7_10);
	-- signal N0_7_11 : std_logic;
	PP376 : and2 port map (X(4), Y(7), N0_7_11);
	-- signal N0_7_12 : std_logic;
	PP377 : and2 port map (X(5), Y(7), N0_7_12);
	-- signal N0_7_13 : std_logic;
	PP378 : and2 port map (X(6), Y(7), N0_7_13);
	-- signal N0_7_14 : std_logic;
	PP379 : and2 port map (X(7), Y(7), N0_7_14);
	-- signal N0_7_15 : std_logic;
	PP380 : and2 port map (X(8), Y(7), N0_7_15);
	-- signal N0_7_16 : std_logic;
	PP381 : and2 port map (X(9), Y(7), N0_7_16);
	-- signal N0_7_17 : std_logic;
	PP382 : and2 port map (X(10), Y(7), N0_7_17);
	-- signal N0_7_18 : std_logic;
	PP383 : and2 port map (X(11), Y(7), N0_7_18);
	-- signal N0_7_19 : std_logic;
	PP384 : and2 port map (X(12), Y(7), N0_7_19);
	-- signal N0_7_20 : std_logic;
	PP385 : and2 port map (X(13), Y(7), N0_7_20);
	-- signal N0_7_21 : std_logic;
	PP386 : and2 port map (X(14), Y(7), N0_7_21);
	-- signal N0_7_22 : std_logic;
	PP387 : and2 port map (X(15), Y(7), N0_7_22);
	-- signal N0_7_23 : std_logic;
	PP388 : and2 port map (X(16), Y(7), N0_7_23);
	-- signal N0_7_24 : std_logic;
	PP389 : and2 port map (X(17), Y(7), N0_7_24);
	-- signal N0_7_25 : std_logic;
	PP390 : and2 port map (X(18), Y(7), N0_7_25);
	-- signal N0_7_26 : std_logic;
	PP391 : and2 port map (X(19), Y(7), N0_7_26);
	-- signal N0_7_27 : std_logic;
	PP392 : and2 port map (X(20), Y(7), N0_7_27);
	-- signal N0_7_28 : std_logic;
	PP393 : and2 port map (X(21), Y(7), N0_7_28);
	-- signal N0_7_29 : std_logic;
	PP394 : and2 port map (X(22), Y(7), N0_7_29);
	-- signal N0_7_30 : std_logic;
	PP395 : and2 port map (X(23), Y(7), N0_7_30);
	-- signal N0_7_31 : std_logic;
	PP396 : and2 port map (X(24), Y(7), N0_7_31);
	-- signal N0_7_32 : std_logic;
	PP397 : and2 port map (X(25), Y(7), N0_7_32);
	-- signal N0_7_33 : std_logic;
	PP398 : and2 port map (X(26), Y(7), N0_7_33);
	-- signal N0_7_34 : std_logic;
	PP399 : and2 port map (X(27), Y(7), N0_7_34);
	-- signal N0_7_35 : std_logic;
	PP400 : and2 port map (X(28), Y(7), N0_7_35);
	-- signal N0_7_36 : std_logic;
	PP401 : and2 port map (X(29), Y(7), N0_7_36);
	-- signal N0_7_37 : std_logic;
	PP402 : and2 port map (X(30), Y(7), N0_7_37);
	-- signal N0_7_38 : std_logic;
	PP403 : and2 port map (X(31), Y(7), N0_7_38);
	-- signal N0_7_39 : std_logic;
	PP404 : and2 port map (X(32), Y(7), N0_7_39);
	-- signal N0_7_40 : std_logic;
	PP405 : and2 port map (X(33), Y(7), N0_7_40);
	-- signal N0_7_41 : std_logic;
	PP406 : and2 port map (X(34), Y(7), N0_7_41);
	-- signal N0_7_42 : std_logic;
	PP407 : and2 port map (X(35), Y(7), N0_7_42);
	-- signal N0_7_43 : std_logic;
	PP408 : and2 port map (X(36), Y(7), N0_7_43);
	-- signal N0_7_44 : std_logic;
	PP409 : and2 port map (X(37), Y(7), N0_7_44);
	-- signal N0_7_45 : std_logic;
	PP410 : and2 port map (X(38), Y(7), N0_7_45);
	-- signal N0_7_46 : std_logic;
	PP411 : and2 port map (X(39), Y(7), N0_7_46);
	-- signal N0_7_47 : std_logic;
	PP412 : and2 port map (X(40), Y(7), N0_7_47);
	-- signal N0_7_48 : std_logic;
	PP413 : and2 port map (X(41), Y(7), N0_7_48);
	-- signal N0_7_49 : std_logic;
	PP414 : and2 port map (X(42), Y(7), N0_7_49);
	-- signal N0_7_50 : std_logic;
	PP415 : and2 port map (X(43), Y(7), N0_7_50);
	-- signal N0_7_51 : std_logic;
	PP416 : and2 port map (X(44), Y(7), N0_7_51);
	-- signal N0_7_52 : std_logic;
	PP417 : and2 port map (X(45), Y(7), N0_7_52);
	-- signal N0_7_53 : std_logic;
	PP418 : and2 port map (X(46), Y(7), N0_7_53);
	-- signal N0_7_54 : std_logic;
	PP419 : and2 port map (X(47), Y(7), N0_7_54);
	-- signal N0_7_55 : std_logic;
	PP420 : and2 port map (X(48), Y(7), N0_7_55);
	-- signal N0_7_56 : std_logic;
	PP421 : and2 port map (X(49), Y(7), N0_7_56);
	-- signal N0_7_57 : std_logic;
	PP422 : and2 port map (X(50), Y(7), N0_7_57);
	-- signal N0_7_58 : std_logic;
	PP423 : and2 port map (X(51), Y(7), N0_7_58);
	-- signal N0_7_59 : std_logic;
	PP424 : and2 port map ('1', Y(7), N0_7_59);
	-- signal N0_8_8 : std_logic;
	PP425 : and2 port map (X(0), Y(8), N0_8_8);
	-- signal N0_8_9 : std_logic;
	PP426 : and2 port map (X(1), Y(8), N0_8_9);
	-- signal N0_8_10 : std_logic;
	PP427 : and2 port map (X(2), Y(8), N0_8_10);
	-- signal N0_8_11 : std_logic;
	PP428 : and2 port map (X(3), Y(8), N0_8_11);
	-- signal N0_8_12 : std_logic;
	PP429 : and2 port map (X(4), Y(8), N0_8_12);
	-- signal N0_8_13 : std_logic;
	PP430 : and2 port map (X(5), Y(8), N0_8_13);
	-- signal N0_8_14 : std_logic;
	PP431 : and2 port map (X(6), Y(8), N0_8_14);
	-- signal N0_8_15 : std_logic;
	PP432 : and2 port map (X(7), Y(8), N0_8_15);
	-- signal N0_8_16 : std_logic;
	PP433 : and2 port map (X(8), Y(8), N0_8_16);
	-- signal N0_8_17 : std_logic;
	PP434 : and2 port map (X(9), Y(8), N0_8_17);
	-- signal N0_8_18 : std_logic;
	PP435 : and2 port map (X(10), Y(8), N0_8_18);
	-- signal N0_8_19 : std_logic;
	PP436 : and2 port map (X(11), Y(8), N0_8_19);
	-- signal N0_8_20 : std_logic;
	PP437 : and2 port map (X(12), Y(8), N0_8_20);
	-- signal N0_8_21 : std_logic;
	PP438 : and2 port map (X(13), Y(8), N0_8_21);
	-- signal N0_8_22 : std_logic;
	PP439 : and2 port map (X(14), Y(8), N0_8_22);
	-- signal N0_8_23 : std_logic;
	PP440 : and2 port map (X(15), Y(8), N0_8_23);
	-- signal N0_8_24 : std_logic;
	PP441 : and2 port map (X(16), Y(8), N0_8_24);
	-- signal N0_8_25 : std_logic;
	PP442 : and2 port map (X(17), Y(8), N0_8_25);
	-- signal N0_8_26 : std_logic;
	PP443 : and2 port map (X(18), Y(8), N0_8_26);
	-- signal N0_8_27 : std_logic;
	PP444 : and2 port map (X(19), Y(8), N0_8_27);
	-- signal N0_8_28 : std_logic;
	PP445 : and2 port map (X(20), Y(8), N0_8_28);
	-- signal N0_8_29 : std_logic;
	PP446 : and2 port map (X(21), Y(8), N0_8_29);
	-- signal N0_8_30 : std_logic;
	PP447 : and2 port map (X(22), Y(8), N0_8_30);
	-- signal N0_8_31 : std_logic;
	PP448 : and2 port map (X(23), Y(8), N0_8_31);
	-- signal N0_8_32 : std_logic;
	PP449 : and2 port map (X(24), Y(8), N0_8_32);
	-- signal N0_8_33 : std_logic;
	PP450 : and2 port map (X(25), Y(8), N0_8_33);
	-- signal N0_8_34 : std_logic;
	PP451 : and2 port map (X(26), Y(8), N0_8_34);
	-- signal N0_8_35 : std_logic;
	PP452 : and2 port map (X(27), Y(8), N0_8_35);
	-- signal N0_8_36 : std_logic;
	PP453 : and2 port map (X(28), Y(8), N0_8_36);
	-- signal N0_8_37 : std_logic;
	PP454 : and2 port map (X(29), Y(8), N0_8_37);
	-- signal N0_8_38 : std_logic;
	PP455 : and2 port map (X(30), Y(8), N0_8_38);
	-- signal N0_8_39 : std_logic;
	PP456 : and2 port map (X(31), Y(8), N0_8_39);
	-- signal N0_8_40 : std_logic;
	PP457 : and2 port map (X(32), Y(8), N0_8_40);
	-- signal N0_8_41 : std_logic;
	PP458 : and2 port map (X(33), Y(8), N0_8_41);
	-- signal N0_8_42 : std_logic;
	PP459 : and2 port map (X(34), Y(8), N0_8_42);
	-- signal N0_8_43 : std_logic;
	PP460 : and2 port map (X(35), Y(8), N0_8_43);
	-- signal N0_8_44 : std_logic;
	PP461 : and2 port map (X(36), Y(8), N0_8_44);
	-- signal N0_8_45 : std_logic;
	PP462 : and2 port map (X(37), Y(8), N0_8_45);
	-- signal N0_8_46 : std_logic;
	PP463 : and2 port map (X(38), Y(8), N0_8_46);
	-- signal N0_8_47 : std_logic;
	PP464 : and2 port map (X(39), Y(8), N0_8_47);
	-- signal N0_8_48 : std_logic;
	PP465 : and2 port map (X(40), Y(8), N0_8_48);
	-- signal N0_8_49 : std_logic;
	PP466 : and2 port map (X(41), Y(8), N0_8_49);
	-- signal N0_8_50 : std_logic;
	PP467 : and2 port map (X(42), Y(8), N0_8_50);
	-- signal N0_8_51 : std_logic;
	PP468 : and2 port map (X(43), Y(8), N0_8_51);
	-- signal N0_8_52 : std_logic;
	PP469 : and2 port map (X(44), Y(8), N0_8_52);
	-- signal N0_8_53 : std_logic;
	PP470 : and2 port map (X(45), Y(8), N0_8_53);
	-- signal N0_8_54 : std_logic;
	PP471 : and2 port map (X(46), Y(8), N0_8_54);
	-- signal N0_8_55 : std_logic;
	PP472 : and2 port map (X(47), Y(8), N0_8_55);
	-- signal N0_8_56 : std_logic;
	PP473 : and2 port map (X(48), Y(8), N0_8_56);
	-- signal N0_8_57 : std_logic;
	PP474 : and2 port map (X(49), Y(8), N0_8_57);
	-- signal N0_8_58 : std_logic;
	PP475 : and2 port map (X(50), Y(8), N0_8_58);
	-- signal N0_8_59 : std_logic;
	PP476 : and2 port map (X(51), Y(8), N0_8_59);
	-- signal N0_8_60 : std_logic;
	PP477 : and2 port map ('1', Y(8), N0_8_60);
	-- signal N0_9_9 : std_logic;
	PP478 : and2 port map (X(0), Y(9), N0_9_9);
	-- signal N0_9_10 : std_logic;
	PP479 : and2 port map (X(1), Y(9), N0_9_10);
	-- signal N0_9_11 : std_logic;
	PP480 : and2 port map (X(2), Y(9), N0_9_11);
	-- signal N0_9_12 : std_logic;
	PP481 : and2 port map (X(3), Y(9), N0_9_12);
	-- signal N0_9_13 : std_logic;
	PP482 : and2 port map (X(4), Y(9), N0_9_13);
	-- signal N0_9_14 : std_logic;
	PP483 : and2 port map (X(5), Y(9), N0_9_14);
	-- signal N0_9_15 : std_logic;
	PP484 : and2 port map (X(6), Y(9), N0_9_15);
	-- signal N0_9_16 : std_logic;
	PP485 : and2 port map (X(7), Y(9), N0_9_16);
	-- signal N0_9_17 : std_logic;
	PP486 : and2 port map (X(8), Y(9), N0_9_17);
	-- signal N0_9_18 : std_logic;
	PP487 : and2 port map (X(9), Y(9), N0_9_18);
	-- signal N0_9_19 : std_logic;
	PP488 : and2 port map (X(10), Y(9), N0_9_19);
	-- signal N0_9_20 : std_logic;
	PP489 : and2 port map (X(11), Y(9), N0_9_20);
	-- signal N0_9_21 : std_logic;
	PP490 : and2 port map (X(12), Y(9), N0_9_21);
	-- signal N0_9_22 : std_logic;
	PP491 : and2 port map (X(13), Y(9), N0_9_22);
	-- signal N0_9_23 : std_logic;
	PP492 : and2 port map (X(14), Y(9), N0_9_23);
	-- signal N0_9_24 : std_logic;
	PP493 : and2 port map (X(15), Y(9), N0_9_24);
	-- signal N0_9_25 : std_logic;
	PP494 : and2 port map (X(16), Y(9), N0_9_25);
	-- signal N0_9_26 : std_logic;
	PP495 : and2 port map (X(17), Y(9), N0_9_26);
	-- signal N0_9_27 : std_logic;
	PP496 : and2 port map (X(18), Y(9), N0_9_27);
	-- signal N0_9_28 : std_logic;
	PP497 : and2 port map (X(19), Y(9), N0_9_28);
	-- signal N0_9_29 : std_logic;
	PP498 : and2 port map (X(20), Y(9), N0_9_29);
	-- signal N0_9_30 : std_logic;
	PP499 : and2 port map (X(21), Y(9), N0_9_30);
	-- signal N0_9_31 : std_logic;
	PP500 : and2 port map (X(22), Y(9), N0_9_31);
	-- signal N0_9_32 : std_logic;
	PP501 : and2 port map (X(23), Y(9), N0_9_32);
	-- signal N0_9_33 : std_logic;
	PP502 : and2 port map (X(24), Y(9), N0_9_33);
	-- signal N0_9_34 : std_logic;
	PP503 : and2 port map (X(25), Y(9), N0_9_34);
	-- signal N0_9_35 : std_logic;
	PP504 : and2 port map (X(26), Y(9), N0_9_35);
	-- signal N0_9_36 : std_logic;
	PP505 : and2 port map (X(27), Y(9), N0_9_36);
	-- signal N0_9_37 : std_logic;
	PP506 : and2 port map (X(28), Y(9), N0_9_37);
	-- signal N0_9_38 : std_logic;
	PP507 : and2 port map (X(29), Y(9), N0_9_38);
	-- signal N0_9_39 : std_logic;
	PP508 : and2 port map (X(30), Y(9), N0_9_39);
	-- signal N0_9_40 : std_logic;
	PP509 : and2 port map (X(31), Y(9), N0_9_40);
	-- signal N0_9_41 : std_logic;
	PP510 : and2 port map (X(32), Y(9), N0_9_41);
	-- signal N0_9_42 : std_logic;
	PP511 : and2 port map (X(33), Y(9), N0_9_42);
	-- signal N0_9_43 : std_logic;
	PP512 : and2 port map (X(34), Y(9), N0_9_43);
	-- signal N0_9_44 : std_logic;
	PP513 : and2 port map (X(35), Y(9), N0_9_44);
	-- signal N0_9_45 : std_logic;
	PP514 : and2 port map (X(36), Y(9), N0_9_45);
	-- signal N0_9_46 : std_logic;
	PP515 : and2 port map (X(37), Y(9), N0_9_46);
	-- signal N0_9_47 : std_logic;
	PP516 : and2 port map (X(38), Y(9), N0_9_47);
	-- signal N0_9_48 : std_logic;
	PP517 : and2 port map (X(39), Y(9), N0_9_48);
	-- signal N0_9_49 : std_logic;
	PP518 : and2 port map (X(40), Y(9), N0_9_49);
	-- signal N0_9_50 : std_logic;
	PP519 : and2 port map (X(41), Y(9), N0_9_50);
	-- signal N0_9_51 : std_logic;
	PP520 : and2 port map (X(42), Y(9), N0_9_51);
	-- signal N0_9_52 : std_logic;
	PP521 : and2 port map (X(43), Y(9), N0_9_52);
	-- signal N0_9_53 : std_logic;
	PP522 : and2 port map (X(44), Y(9), N0_9_53);
	-- signal N0_9_54 : std_logic;
	PP523 : and2 port map (X(45), Y(9), N0_9_54);
	-- signal N0_9_55 : std_logic;
	PP524 : and2 port map (X(46), Y(9), N0_9_55);
	-- signal N0_9_56 : std_logic;
	PP525 : and2 port map (X(47), Y(9), N0_9_56);
	-- signal N0_9_57 : std_logic;
	PP526 : and2 port map (X(48), Y(9), N0_9_57);
	-- signal N0_9_58 : std_logic;
	PP527 : and2 port map (X(49), Y(9), N0_9_58);
	-- signal N0_9_59 : std_logic;
	PP528 : and2 port map (X(50), Y(9), N0_9_59);
	-- signal N0_9_60 : std_logic;
	PP529 : and2 port map (X(51), Y(9), N0_9_60);
	-- signal N0_9_61 : std_logic;
	PP530 : and2 port map ('1', Y(9), N0_9_61);
	-- signal N0_10_10 : std_logic;
	PP531 : and2 port map (X(0), Y(10), N0_10_10);
	-- signal N0_10_11 : std_logic;
	PP532 : and2 port map (X(1), Y(10), N0_10_11);
	-- signal N0_10_12 : std_logic;
	PP533 : and2 port map (X(2), Y(10), N0_10_12);
	-- signal N0_10_13 : std_logic;
	PP534 : and2 port map (X(3), Y(10), N0_10_13);
	-- signal N0_10_14 : std_logic;
	PP535 : and2 port map (X(4), Y(10), N0_10_14);
	-- signal N0_10_15 : std_logic;
	PP536 : and2 port map (X(5), Y(10), N0_10_15);
	-- signal N0_10_16 : std_logic;
	PP537 : and2 port map (X(6), Y(10), N0_10_16);
	-- signal N0_10_17 : std_logic;
	PP538 : and2 port map (X(7), Y(10), N0_10_17);
	-- signal N0_10_18 : std_logic;
	PP539 : and2 port map (X(8), Y(10), N0_10_18);
	-- signal N0_10_19 : std_logic;
	PP540 : and2 port map (X(9), Y(10), N0_10_19);
	-- signal N0_10_20 : std_logic;
	PP541 : and2 port map (X(10), Y(10), N0_10_20);
	-- signal N0_10_21 : std_logic;
	PP542 : and2 port map (X(11), Y(10), N0_10_21);
	-- signal N0_10_22 : std_logic;
	PP543 : and2 port map (X(12), Y(10), N0_10_22);
	-- signal N0_10_23 : std_logic;
	PP544 : and2 port map (X(13), Y(10), N0_10_23);
	-- signal N0_10_24 : std_logic;
	PP545 : and2 port map (X(14), Y(10), N0_10_24);
	-- signal N0_10_25 : std_logic;
	PP546 : and2 port map (X(15), Y(10), N0_10_25);
	-- signal N0_10_26 : std_logic;
	PP547 : and2 port map (X(16), Y(10), N0_10_26);
	-- signal N0_10_27 : std_logic;
	PP548 : and2 port map (X(17), Y(10), N0_10_27);
	-- signal N0_10_28 : std_logic;
	PP549 : and2 port map (X(18), Y(10), N0_10_28);
	-- signal N0_10_29 : std_logic;
	PP550 : and2 port map (X(19), Y(10), N0_10_29);
	-- signal N0_10_30 : std_logic;
	PP551 : and2 port map (X(20), Y(10), N0_10_30);
	-- signal N0_10_31 : std_logic;
	PP552 : and2 port map (X(21), Y(10), N0_10_31);
	-- signal N0_10_32 : std_logic;
	PP553 : and2 port map (X(22), Y(10), N0_10_32);
	-- signal N0_10_33 : std_logic;
	PP554 : and2 port map (X(23), Y(10), N0_10_33);
	-- signal N0_10_34 : std_logic;
	PP555 : and2 port map (X(24), Y(10), N0_10_34);
	-- signal N0_10_35 : std_logic;
	PP556 : and2 port map (X(25), Y(10), N0_10_35);
	-- signal N0_10_36 : std_logic;
	PP557 : and2 port map (X(26), Y(10), N0_10_36);
	-- signal N0_10_37 : std_logic;
	PP558 : and2 port map (X(27), Y(10), N0_10_37);
	-- signal N0_10_38 : std_logic;
	PP559 : and2 port map (X(28), Y(10), N0_10_38);
	-- signal N0_10_39 : std_logic;
	PP560 : and2 port map (X(29), Y(10), N0_10_39);
	-- signal N0_10_40 : std_logic;
	PP561 : and2 port map (X(30), Y(10), N0_10_40);
	-- signal N0_10_41 : std_logic;
	PP562 : and2 port map (X(31), Y(10), N0_10_41);
	-- signal N0_10_42 : std_logic;
	PP563 : and2 port map (X(32), Y(10), N0_10_42);
	-- signal N0_10_43 : std_logic;
	PP564 : and2 port map (X(33), Y(10), N0_10_43);
	-- signal N0_10_44 : std_logic;
	PP565 : and2 port map (X(34), Y(10), N0_10_44);
	-- signal N0_10_45 : std_logic;
	PP566 : and2 port map (X(35), Y(10), N0_10_45);
	-- signal N0_10_46 : std_logic;
	PP567 : and2 port map (X(36), Y(10), N0_10_46);
	-- signal N0_10_47 : std_logic;
	PP568 : and2 port map (X(37), Y(10), N0_10_47);
	-- signal N0_10_48 : std_logic;
	PP569 : and2 port map (X(38), Y(10), N0_10_48);
	-- signal N0_10_49 : std_logic;
	PP570 : and2 port map (X(39), Y(10), N0_10_49);
	-- signal N0_10_50 : std_logic;
	PP571 : and2 port map (X(40), Y(10), N0_10_50);
	-- signal N0_10_51 : std_logic;
	PP572 : and2 port map (X(41), Y(10), N0_10_51);
	-- signal N0_10_52 : std_logic;
	PP573 : and2 port map (X(42), Y(10), N0_10_52);
	-- signal N0_10_53 : std_logic;
	PP574 : and2 port map (X(43), Y(10), N0_10_53);
	-- signal N0_10_54 : std_logic;
	PP575 : and2 port map (X(44), Y(10), N0_10_54);
	-- signal N0_10_55 : std_logic;
	PP576 : and2 port map (X(45), Y(10), N0_10_55);
	-- signal N0_10_56 : std_logic;
	PP577 : and2 port map (X(46), Y(10), N0_10_56);
	-- signal N0_10_57 : std_logic;
	PP578 : and2 port map (X(47), Y(10), N0_10_57);
	-- signal N0_10_58 : std_logic;
	PP579 : and2 port map (X(48), Y(10), N0_10_58);
	-- signal N0_10_59 : std_logic;
	PP580 : and2 port map (X(49), Y(10), N0_10_59);
	-- signal N0_10_60 : std_logic;
	PP581 : and2 port map (X(50), Y(10), N0_10_60);
	-- signal N0_10_61 : std_logic;
	PP582 : and2 port map (X(51), Y(10), N0_10_61);
	-- signal N0_10_62 : std_logic;
	PP583 : and2 port map ('1', Y(10), N0_10_62);
	-- signal N0_11_11 : std_logic;
	PP584 : and2 port map (X(0), Y(11), N0_11_11);
	-- signal N0_11_12 : std_logic;
	PP585 : and2 port map (X(1), Y(11), N0_11_12);
	-- signal N0_11_13 : std_logic;
	PP586 : and2 port map (X(2), Y(11), N0_11_13);
	-- signal N0_11_14 : std_logic;
	PP587 : and2 port map (X(3), Y(11), N0_11_14);
	-- signal N0_11_15 : std_logic;
	PP588 : and2 port map (X(4), Y(11), N0_11_15);
	-- signal N0_11_16 : std_logic;
	PP589 : and2 port map (X(5), Y(11), N0_11_16);
	-- signal N0_11_17 : std_logic;
	PP590 : and2 port map (X(6), Y(11), N0_11_17);
	-- signal N0_11_18 : std_logic;
	PP591 : and2 port map (X(7), Y(11), N0_11_18);
	-- signal N0_11_19 : std_logic;
	PP592 : and2 port map (X(8), Y(11), N0_11_19);
	-- signal N0_11_20 : std_logic;
	PP593 : and2 port map (X(9), Y(11), N0_11_20);
	-- signal N0_11_21 : std_logic;
	PP594 : and2 port map (X(10), Y(11), N0_11_21);
	-- signal N0_11_22 : std_logic;
	PP595 : and2 port map (X(11), Y(11), N0_11_22);
	-- signal N0_11_23 : std_logic;
	PP596 : and2 port map (X(12), Y(11), N0_11_23);
	-- signal N0_11_24 : std_logic;
	PP597 : and2 port map (X(13), Y(11), N0_11_24);
	-- signal N0_11_25 : std_logic;
	PP598 : and2 port map (X(14), Y(11), N0_11_25);
	-- signal N0_11_26 : std_logic;
	PP599 : and2 port map (X(15), Y(11), N0_11_26);
	-- signal N0_11_27 : std_logic;
	PP600 : and2 port map (X(16), Y(11), N0_11_27);
	-- signal N0_11_28 : std_logic;
	PP601 : and2 port map (X(17), Y(11), N0_11_28);
	-- signal N0_11_29 : std_logic;
	PP602 : and2 port map (X(18), Y(11), N0_11_29);
	-- signal N0_11_30 : std_logic;
	PP603 : and2 port map (X(19), Y(11), N0_11_30);
	-- signal N0_11_31 : std_logic;
	PP604 : and2 port map (X(20), Y(11), N0_11_31);
	-- signal N0_11_32 : std_logic;
	PP605 : and2 port map (X(21), Y(11), N0_11_32);
	-- signal N0_11_33 : std_logic;
	PP606 : and2 port map (X(22), Y(11), N0_11_33);
	-- signal N0_11_34 : std_logic;
	PP607 : and2 port map (X(23), Y(11), N0_11_34);
	-- signal N0_11_35 : std_logic;
	PP608 : and2 port map (X(24), Y(11), N0_11_35);
	-- signal N0_11_36 : std_logic;
	PP609 : and2 port map (X(25), Y(11), N0_11_36);
	-- signal N0_11_37 : std_logic;
	PP610 : and2 port map (X(26), Y(11), N0_11_37);
	-- signal N0_11_38 : std_logic;
	PP611 : and2 port map (X(27), Y(11), N0_11_38);
	-- signal N0_11_39 : std_logic;
	PP612 : and2 port map (X(28), Y(11), N0_11_39);
	-- signal N0_11_40 : std_logic;
	PP613 : and2 port map (X(29), Y(11), N0_11_40);
	-- signal N0_11_41 : std_logic;
	PP614 : and2 port map (X(30), Y(11), N0_11_41);
	-- signal N0_11_42 : std_logic;
	PP615 : and2 port map (X(31), Y(11), N0_11_42);
	-- signal N0_11_43 : std_logic;
	PP616 : and2 port map (X(32), Y(11), N0_11_43);
	-- signal N0_11_44 : std_logic;
	PP617 : and2 port map (X(33), Y(11), N0_11_44);
	-- signal N0_11_45 : std_logic;
	PP618 : and2 port map (X(34), Y(11), N0_11_45);
	-- signal N0_11_46 : std_logic;
	PP619 : and2 port map (X(35), Y(11), N0_11_46);
	-- signal N0_11_47 : std_logic;
	PP620 : and2 port map (X(36), Y(11), N0_11_47);
	-- signal N0_11_48 : std_logic;
	PP621 : and2 port map (X(37), Y(11), N0_11_48);
	-- signal N0_11_49 : std_logic;
	PP622 : and2 port map (X(38), Y(11), N0_11_49);
	-- signal N0_11_50 : std_logic;
	PP623 : and2 port map (X(39), Y(11), N0_11_50);
	-- signal N0_11_51 : std_logic;
	PP624 : and2 port map (X(40), Y(11), N0_11_51);
	-- signal N0_11_52 : std_logic;
	PP625 : and2 port map (X(41), Y(11), N0_11_52);
	-- signal N0_11_53 : std_logic;
	PP626 : and2 port map (X(42), Y(11), N0_11_53);
	-- signal N0_11_54 : std_logic;
	PP627 : and2 port map (X(43), Y(11), N0_11_54);
	-- signal N0_11_55 : std_logic;
	PP628 : and2 port map (X(44), Y(11), N0_11_55);
	-- signal N0_11_56 : std_logic;
	PP629 : and2 port map (X(45), Y(11), N0_11_56);
	-- signal N0_11_57 : std_logic;
	PP630 : and2 port map (X(46), Y(11), N0_11_57);
	-- signal N0_11_58 : std_logic;
	PP631 : and2 port map (X(47), Y(11), N0_11_58);
	-- signal N0_11_59 : std_logic;
	PP632 : and2 port map (X(48), Y(11), N0_11_59);
	-- signal N0_11_60 : std_logic;
	PP633 : and2 port map (X(49), Y(11), N0_11_60);
	-- signal N0_11_61 : std_logic;
	PP634 : and2 port map (X(50), Y(11), N0_11_61);
	-- signal N0_11_62 : std_logic;
	PP635 : and2 port map (X(51), Y(11), N0_11_62);
	-- signal N0_11_63 : std_logic;
	PP636 : and2 port map ('1', Y(11), N0_11_63);
	-- signal N0_12_12 : std_logic;
	PP637 : and2 port map (X(0), Y(12), N0_12_12);
	-- signal N0_12_13 : std_logic;
	PP638 : and2 port map (X(1), Y(12), N0_12_13);
	-- signal N0_12_14 : std_logic;
	PP639 : and2 port map (X(2), Y(12), N0_12_14);
	-- signal N0_12_15 : std_logic;
	PP640 : and2 port map (X(3), Y(12), N0_12_15);
	-- signal N0_12_16 : std_logic;
	PP641 : and2 port map (X(4), Y(12), N0_12_16);
	-- signal N0_12_17 : std_logic;
	PP642 : and2 port map (X(5), Y(12), N0_12_17);
	-- signal N0_12_18 : std_logic;
	PP643 : and2 port map (X(6), Y(12), N0_12_18);
	-- signal N0_12_19 : std_logic;
	PP644 : and2 port map (X(7), Y(12), N0_12_19);
	-- signal N0_12_20 : std_logic;
	PP645 : and2 port map (X(8), Y(12), N0_12_20);
	-- signal N0_12_21 : std_logic;
	PP646 : and2 port map (X(9), Y(12), N0_12_21);
	-- signal N0_12_22 : std_logic;
	PP647 : and2 port map (X(10), Y(12), N0_12_22);
	-- signal N0_12_23 : std_logic;
	PP648 : and2 port map (X(11), Y(12), N0_12_23);
	-- signal N0_12_24 : std_logic;
	PP649 : and2 port map (X(12), Y(12), N0_12_24);
	-- signal N0_12_25 : std_logic;
	PP650 : and2 port map (X(13), Y(12), N0_12_25);
	-- signal N0_12_26 : std_logic;
	PP651 : and2 port map (X(14), Y(12), N0_12_26);
	-- signal N0_12_27 : std_logic;
	PP652 : and2 port map (X(15), Y(12), N0_12_27);
	-- signal N0_12_28 : std_logic;
	PP653 : and2 port map (X(16), Y(12), N0_12_28);
	-- signal N0_12_29 : std_logic;
	PP654 : and2 port map (X(17), Y(12), N0_12_29);
	-- signal N0_12_30 : std_logic;
	PP655 : and2 port map (X(18), Y(12), N0_12_30);
	-- signal N0_12_31 : std_logic;
	PP656 : and2 port map (X(19), Y(12), N0_12_31);
	-- signal N0_12_32 : std_logic;
	PP657 : and2 port map (X(20), Y(12), N0_12_32);
	-- signal N0_12_33 : std_logic;
	PP658 : and2 port map (X(21), Y(12), N0_12_33);
	-- signal N0_12_34 : std_logic;
	PP659 : and2 port map (X(22), Y(12), N0_12_34);
	-- signal N0_12_35 : std_logic;
	PP660 : and2 port map (X(23), Y(12), N0_12_35);
	-- signal N0_12_36 : std_logic;
	PP661 : and2 port map (X(24), Y(12), N0_12_36);
	-- signal N0_12_37 : std_logic;
	PP662 : and2 port map (X(25), Y(12), N0_12_37);
	-- signal N0_12_38 : std_logic;
	PP663 : and2 port map (X(26), Y(12), N0_12_38);
	-- signal N0_12_39 : std_logic;
	PP664 : and2 port map (X(27), Y(12), N0_12_39);
	-- signal N0_12_40 : std_logic;
	PP665 : and2 port map (X(28), Y(12), N0_12_40);
	-- signal N0_12_41 : std_logic;
	PP666 : and2 port map (X(29), Y(12), N0_12_41);
	-- signal N0_12_42 : std_logic;
	PP667 : and2 port map (X(30), Y(12), N0_12_42);
	-- signal N0_12_43 : std_logic;
	PP668 : and2 port map (X(31), Y(12), N0_12_43);
	-- signal N0_12_44 : std_logic;
	PP669 : and2 port map (X(32), Y(12), N0_12_44);
	-- signal N0_12_45 : std_logic;
	PP670 : and2 port map (X(33), Y(12), N0_12_45);
	-- signal N0_12_46 : std_logic;
	PP671 : and2 port map (X(34), Y(12), N0_12_46);
	-- signal N0_12_47 : std_logic;
	PP672 : and2 port map (X(35), Y(12), N0_12_47);
	-- signal N0_12_48 : std_logic;
	PP673 : and2 port map (X(36), Y(12), N0_12_48);
	-- signal N0_12_49 : std_logic;
	PP674 : and2 port map (X(37), Y(12), N0_12_49);
	-- signal N0_12_50 : std_logic;
	PP675 : and2 port map (X(38), Y(12), N0_12_50);
	-- signal N0_12_51 : std_logic;
	PP676 : and2 port map (X(39), Y(12), N0_12_51);
	-- signal N0_12_52 : std_logic;
	PP677 : and2 port map (X(40), Y(12), N0_12_52);
	-- signal N0_12_53 : std_logic;
	PP678 : and2 port map (X(41), Y(12), N0_12_53);
	-- signal N0_12_54 : std_logic;
	PP679 : and2 port map (X(42), Y(12), N0_12_54);
	-- signal N0_12_55 : std_logic;
	PP680 : and2 port map (X(43), Y(12), N0_12_55);
	-- signal N0_12_56 : std_logic;
	PP681 : and2 port map (X(44), Y(12), N0_12_56);
	-- signal N0_12_57 : std_logic;
	PP682 : and2 port map (X(45), Y(12), N0_12_57);
	-- signal N0_12_58 : std_logic;
	PP683 : and2 port map (X(46), Y(12), N0_12_58);
	-- signal N0_12_59 : std_logic;
	PP684 : and2 port map (X(47), Y(12), N0_12_59);
	-- signal N0_12_60 : std_logic;
	PP685 : and2 port map (X(48), Y(12), N0_12_60);
	-- signal N0_12_61 : std_logic;
	PP686 : and2 port map (X(49), Y(12), N0_12_61);
	-- signal N0_12_62 : std_logic;
	PP687 : and2 port map (X(50), Y(12), N0_12_62);
	-- signal N0_12_63 : std_logic;
	PP688 : and2 port map (X(51), Y(12), N0_12_63);
	-- signal N0_12_64 : std_logic;
	PP689 : and2 port map ('1', Y(12), N0_12_64);
	-- signal N0_13_13 : std_logic;
	PP690 : and2 port map (X(0), Y(13), N0_13_13);
	-- signal N0_13_14 : std_logic;
	PP691 : and2 port map (X(1), Y(13), N0_13_14);
	-- signal N0_13_15 : std_logic;
	PP692 : and2 port map (X(2), Y(13), N0_13_15);
	-- signal N0_13_16 : std_logic;
	PP693 : and2 port map (X(3), Y(13), N0_13_16);
	-- signal N0_13_17 : std_logic;
	PP694 : and2 port map (X(4), Y(13), N0_13_17);
	-- signal N0_13_18 : std_logic;
	PP695 : and2 port map (X(5), Y(13), N0_13_18);
	-- signal N0_13_19 : std_logic;
	PP696 : and2 port map (X(6), Y(13), N0_13_19);
	-- signal N0_13_20 : std_logic;
	PP697 : and2 port map (X(7), Y(13), N0_13_20);
	-- signal N0_13_21 : std_logic;
	PP698 : and2 port map (X(8), Y(13), N0_13_21);
	-- signal N0_13_22 : std_logic;
	PP699 : and2 port map (X(9), Y(13), N0_13_22);
	-- signal N0_13_23 : std_logic;
	PP700 : and2 port map (X(10), Y(13), N0_13_23);
	-- signal N0_13_24 : std_logic;
	PP701 : and2 port map (X(11), Y(13), N0_13_24);
	-- signal N0_13_25 : std_logic;
	PP702 : and2 port map (X(12), Y(13), N0_13_25);
	-- signal N0_13_26 : std_logic;
	PP703 : and2 port map (X(13), Y(13), N0_13_26);
	-- signal N0_13_27 : std_logic;
	PP704 : and2 port map (X(14), Y(13), N0_13_27);
	-- signal N0_13_28 : std_logic;
	PP705 : and2 port map (X(15), Y(13), N0_13_28);
	-- signal N0_13_29 : std_logic;
	PP706 : and2 port map (X(16), Y(13), N0_13_29);
	-- signal N0_13_30 : std_logic;
	PP707 : and2 port map (X(17), Y(13), N0_13_30);
	-- signal N0_13_31 : std_logic;
	PP708 : and2 port map (X(18), Y(13), N0_13_31);
	-- signal N0_13_32 : std_logic;
	PP709 : and2 port map (X(19), Y(13), N0_13_32);
	-- signal N0_13_33 : std_logic;
	PP710 : and2 port map (X(20), Y(13), N0_13_33);
	-- signal N0_13_34 : std_logic;
	PP711 : and2 port map (X(21), Y(13), N0_13_34);
	-- signal N0_13_35 : std_logic;
	PP712 : and2 port map (X(22), Y(13), N0_13_35);
	-- signal N0_13_36 : std_logic;
	PP713 : and2 port map (X(23), Y(13), N0_13_36);
	-- signal N0_13_37 : std_logic;
	PP714 : and2 port map (X(24), Y(13), N0_13_37);
	-- signal N0_13_38 : std_logic;
	PP715 : and2 port map (X(25), Y(13), N0_13_38);
	-- signal N0_13_39 : std_logic;
	PP716 : and2 port map (X(26), Y(13), N0_13_39);
	-- signal N0_13_40 : std_logic;
	PP717 : and2 port map (X(27), Y(13), N0_13_40);
	-- signal N0_13_41 : std_logic;
	PP718 : and2 port map (X(28), Y(13), N0_13_41);
	-- signal N0_13_42 : std_logic;
	PP719 : and2 port map (X(29), Y(13), N0_13_42);
	-- signal N0_13_43 : std_logic;
	PP720 : and2 port map (X(30), Y(13), N0_13_43);
	-- signal N0_13_44 : std_logic;
	PP721 : and2 port map (X(31), Y(13), N0_13_44);
	-- signal N0_13_45 : std_logic;
	PP722 : and2 port map (X(32), Y(13), N0_13_45);
	-- signal N0_13_46 : std_logic;
	PP723 : and2 port map (X(33), Y(13), N0_13_46);
	-- signal N0_13_47 : std_logic;
	PP724 : and2 port map (X(34), Y(13), N0_13_47);
	-- signal N0_13_48 : std_logic;
	PP725 : and2 port map (X(35), Y(13), N0_13_48);
	-- signal N0_13_49 : std_logic;
	PP726 : and2 port map (X(36), Y(13), N0_13_49);
	-- signal N0_13_50 : std_logic;
	PP727 : and2 port map (X(37), Y(13), N0_13_50);
	-- signal N0_13_51 : std_logic;
	PP728 : and2 port map (X(38), Y(13), N0_13_51);
	-- signal N0_13_52 : std_logic;
	PP729 : and2 port map (X(39), Y(13), N0_13_52);
	-- signal N0_13_53 : std_logic;
	PP730 : and2 port map (X(40), Y(13), N0_13_53);
	-- signal N0_13_54 : std_logic;
	PP731 : and2 port map (X(41), Y(13), N0_13_54);
	-- signal N0_13_55 : std_logic;
	PP732 : and2 port map (X(42), Y(13), N0_13_55);
	-- signal N0_13_56 : std_logic;
	PP733 : and2 port map (X(43), Y(13), N0_13_56);
	-- signal N0_13_57 : std_logic;
	PP734 : and2 port map (X(44), Y(13), N0_13_57);
	-- signal N0_13_58 : std_logic;
	PP735 : and2 port map (X(45), Y(13), N0_13_58);
	-- signal N0_13_59 : std_logic;
	PP736 : and2 port map (X(46), Y(13), N0_13_59);
	-- signal N0_13_60 : std_logic;
	PP737 : and2 port map (X(47), Y(13), N0_13_60);
	-- signal N0_13_61 : std_logic;
	PP738 : and2 port map (X(48), Y(13), N0_13_61);
	-- signal N0_13_62 : std_logic;
	PP739 : and2 port map (X(49), Y(13), N0_13_62);
	-- signal N0_13_63 : std_logic;
	PP740 : and2 port map (X(50), Y(13), N0_13_63);
	-- signal N0_13_64 : std_logic;
	PP741 : and2 port map (X(51), Y(13), N0_13_64);
	-- signal N0_13_65 : std_logic;
	PP742 : and2 port map ('1', Y(13), N0_13_65);
	-- signal N0_14_14 : std_logic;
	PP743 : and2 port map (X(0), Y(14), N0_14_14);
	-- signal N0_14_15 : std_logic;
	PP744 : and2 port map (X(1), Y(14), N0_14_15);
	-- signal N0_14_16 : std_logic;
	PP745 : and2 port map (X(2), Y(14), N0_14_16);
	-- signal N0_14_17 : std_logic;
	PP746 : and2 port map (X(3), Y(14), N0_14_17);
	-- signal N0_14_18 : std_logic;
	PP747 : and2 port map (X(4), Y(14), N0_14_18);
	-- signal N0_14_19 : std_logic;
	PP748 : and2 port map (X(5), Y(14), N0_14_19);
	-- signal N0_14_20 : std_logic;
	PP749 : and2 port map (X(6), Y(14), N0_14_20);
	-- signal N0_14_21 : std_logic;
	PP750 : and2 port map (X(7), Y(14), N0_14_21);
	-- signal N0_14_22 : std_logic;
	PP751 : and2 port map (X(8), Y(14), N0_14_22);
	-- signal N0_14_23 : std_logic;
	PP752 : and2 port map (X(9), Y(14), N0_14_23);
	-- signal N0_14_24 : std_logic;
	PP753 : and2 port map (X(10), Y(14), N0_14_24);
	-- signal N0_14_25 : std_logic;
	PP754 : and2 port map (X(11), Y(14), N0_14_25);
	-- signal N0_14_26 : std_logic;
	PP755 : and2 port map (X(12), Y(14), N0_14_26);
	-- signal N0_14_27 : std_logic;
	PP756 : and2 port map (X(13), Y(14), N0_14_27);
	-- signal N0_14_28 : std_logic;
	PP757 : and2 port map (X(14), Y(14), N0_14_28);
	-- signal N0_14_29 : std_logic;
	PP758 : and2 port map (X(15), Y(14), N0_14_29);
	-- signal N0_14_30 : std_logic;
	PP759 : and2 port map (X(16), Y(14), N0_14_30);
	-- signal N0_14_31 : std_logic;
	PP760 : and2 port map (X(17), Y(14), N0_14_31);
	-- signal N0_14_32 : std_logic;
	PP761 : and2 port map (X(18), Y(14), N0_14_32);
	-- signal N0_14_33 : std_logic;
	PP762 : and2 port map (X(19), Y(14), N0_14_33);
	-- signal N0_14_34 : std_logic;
	PP763 : and2 port map (X(20), Y(14), N0_14_34);
	-- signal N0_14_35 : std_logic;
	PP764 : and2 port map (X(21), Y(14), N0_14_35);
	-- signal N0_14_36 : std_logic;
	PP765 : and2 port map (X(22), Y(14), N0_14_36);
	-- signal N0_14_37 : std_logic;
	PP766 : and2 port map (X(23), Y(14), N0_14_37);
	-- signal N0_14_38 : std_logic;
	PP767 : and2 port map (X(24), Y(14), N0_14_38);
	-- signal N0_14_39 : std_logic;
	PP768 : and2 port map (X(25), Y(14), N0_14_39);
	-- signal N0_14_40 : std_logic;
	PP769 : and2 port map (X(26), Y(14), N0_14_40);
	-- signal N0_14_41 : std_logic;
	PP770 : and2 port map (X(27), Y(14), N0_14_41);
	-- signal N0_14_42 : std_logic;
	PP771 : and2 port map (X(28), Y(14), N0_14_42);
	-- signal N0_14_43 : std_logic;
	PP772 : and2 port map (X(29), Y(14), N0_14_43);
	-- signal N0_14_44 : std_logic;
	PP773 : and2 port map (X(30), Y(14), N0_14_44);
	-- signal N0_14_45 : std_logic;
	PP774 : and2 port map (X(31), Y(14), N0_14_45);
	-- signal N0_14_46 : std_logic;
	PP775 : and2 port map (X(32), Y(14), N0_14_46);
	-- signal N0_14_47 : std_logic;
	PP776 : and2 port map (X(33), Y(14), N0_14_47);
	-- signal N0_14_48 : std_logic;
	PP777 : and2 port map (X(34), Y(14), N0_14_48);
	-- signal N0_14_49 : std_logic;
	PP778 : and2 port map (X(35), Y(14), N0_14_49);
	-- signal N0_14_50 : std_logic;
	PP779 : and2 port map (X(36), Y(14), N0_14_50);
	-- signal N0_14_51 : std_logic;
	PP780 : and2 port map (X(37), Y(14), N0_14_51);
	-- signal N0_14_52 : std_logic;
	PP781 : and2 port map (X(38), Y(14), N0_14_52);
	-- signal N0_14_53 : std_logic;
	PP782 : and2 port map (X(39), Y(14), N0_14_53);
	-- signal N0_14_54 : std_logic;
	PP783 : and2 port map (X(40), Y(14), N0_14_54);
	-- signal N0_14_55 : std_logic;
	PP784 : and2 port map (X(41), Y(14), N0_14_55);
	-- signal N0_14_56 : std_logic;
	PP785 : and2 port map (X(42), Y(14), N0_14_56);
	-- signal N0_14_57 : std_logic;
	PP786 : and2 port map (X(43), Y(14), N0_14_57);
	-- signal N0_14_58 : std_logic;
	PP787 : and2 port map (X(44), Y(14), N0_14_58);
	-- signal N0_14_59 : std_logic;
	PP788 : and2 port map (X(45), Y(14), N0_14_59);
	-- signal N0_14_60 : std_logic;
	PP789 : and2 port map (X(46), Y(14), N0_14_60);
	-- signal N0_14_61 : std_logic;
	PP790 : and2 port map (X(47), Y(14), N0_14_61);
	-- signal N0_14_62 : std_logic;
	PP791 : and2 port map (X(48), Y(14), N0_14_62);
	-- signal N0_14_63 : std_logic;
	PP792 : and2 port map (X(49), Y(14), N0_14_63);
	-- signal N0_14_64 : std_logic;
	PP793 : and2 port map (X(50), Y(14), N0_14_64);
	-- signal N0_14_65 : std_logic;
	PP794 : and2 port map (X(51), Y(14), N0_14_65);
	-- signal N0_14_66 : std_logic;
	PP795 : and2 port map ('1', Y(14), N0_14_66);
	-- signal N0_15_15 : std_logic;
	PP796 : and2 port map (X(0), Y(15), N0_15_15);
	-- signal N0_15_16 : std_logic;
	PP797 : and2 port map (X(1), Y(15), N0_15_16);
	-- signal N0_15_17 : std_logic;
	PP798 : and2 port map (X(2), Y(15), N0_15_17);
	-- signal N0_15_18 : std_logic;
	PP799 : and2 port map (X(3), Y(15), N0_15_18);
	-- signal N0_15_19 : std_logic;
	PP800 : and2 port map (X(4), Y(15), N0_15_19);
	-- signal N0_15_20 : std_logic;
	PP801 : and2 port map (X(5), Y(15), N0_15_20);
	-- signal N0_15_21 : std_logic;
	PP802 : and2 port map (X(6), Y(15), N0_15_21);
	-- signal N0_15_22 : std_logic;
	PP803 : and2 port map (X(7), Y(15), N0_15_22);
	-- signal N0_15_23 : std_logic;
	PP804 : and2 port map (X(8), Y(15), N0_15_23);
	-- signal N0_15_24 : std_logic;
	PP805 : and2 port map (X(9), Y(15), N0_15_24);
	-- signal N0_15_25 : std_logic;
	PP806 : and2 port map (X(10), Y(15), N0_15_25);
	-- signal N0_15_26 : std_logic;
	PP807 : and2 port map (X(11), Y(15), N0_15_26);
	-- signal N0_15_27 : std_logic;
	PP808 : and2 port map (X(12), Y(15), N0_15_27);
	-- signal N0_15_28 : std_logic;
	PP809 : and2 port map (X(13), Y(15), N0_15_28);
	-- signal N0_15_29 : std_logic;
	PP810 : and2 port map (X(14), Y(15), N0_15_29);
	-- signal N0_15_30 : std_logic;
	PP811 : and2 port map (X(15), Y(15), N0_15_30);
	-- signal N0_15_31 : std_logic;
	PP812 : and2 port map (X(16), Y(15), N0_15_31);
	-- signal N0_15_32 : std_logic;
	PP813 : and2 port map (X(17), Y(15), N0_15_32);
	-- signal N0_15_33 : std_logic;
	PP814 : and2 port map (X(18), Y(15), N0_15_33);
	-- signal N0_15_34 : std_logic;
	PP815 : and2 port map (X(19), Y(15), N0_15_34);
	-- signal N0_15_35 : std_logic;
	PP816 : and2 port map (X(20), Y(15), N0_15_35);
	-- signal N0_15_36 : std_logic;
	PP817 : and2 port map (X(21), Y(15), N0_15_36);
	-- signal N0_15_37 : std_logic;
	PP818 : and2 port map (X(22), Y(15), N0_15_37);
	-- signal N0_15_38 : std_logic;
	PP819 : and2 port map (X(23), Y(15), N0_15_38);
	-- signal N0_15_39 : std_logic;
	PP820 : and2 port map (X(24), Y(15), N0_15_39);
	-- signal N0_15_40 : std_logic;
	PP821 : and2 port map (X(25), Y(15), N0_15_40);
	-- signal N0_15_41 : std_logic;
	PP822 : and2 port map (X(26), Y(15), N0_15_41);
	-- signal N0_15_42 : std_logic;
	PP823 : and2 port map (X(27), Y(15), N0_15_42);
	-- signal N0_15_43 : std_logic;
	PP824 : and2 port map (X(28), Y(15), N0_15_43);
	-- signal N0_15_44 : std_logic;
	PP825 : and2 port map (X(29), Y(15), N0_15_44);
	-- signal N0_15_45 : std_logic;
	PP826 : and2 port map (X(30), Y(15), N0_15_45);
	-- signal N0_15_46 : std_logic;
	PP827 : and2 port map (X(31), Y(15), N0_15_46);
	-- signal N0_15_47 : std_logic;
	PP828 : and2 port map (X(32), Y(15), N0_15_47);
	-- signal N0_15_48 : std_logic;
	PP829 : and2 port map (X(33), Y(15), N0_15_48);
	-- signal N0_15_49 : std_logic;
	PP830 : and2 port map (X(34), Y(15), N0_15_49);
	-- signal N0_15_50 : std_logic;
	PP831 : and2 port map (X(35), Y(15), N0_15_50);
	-- signal N0_15_51 : std_logic;
	PP832 : and2 port map (X(36), Y(15), N0_15_51);
	-- signal N0_15_52 : std_logic;
	PP833 : and2 port map (X(37), Y(15), N0_15_52);
	-- signal N0_15_53 : std_logic;
	PP834 : and2 port map (X(38), Y(15), N0_15_53);
	-- signal N0_15_54 : std_logic;
	PP835 : and2 port map (X(39), Y(15), N0_15_54);
	-- signal N0_15_55 : std_logic;
	PP836 : and2 port map (X(40), Y(15), N0_15_55);
	-- signal N0_15_56 : std_logic;
	PP837 : and2 port map (X(41), Y(15), N0_15_56);
	-- signal N0_15_57 : std_logic;
	PP838 : and2 port map (X(42), Y(15), N0_15_57);
	-- signal N0_15_58 : std_logic;
	PP839 : and2 port map (X(43), Y(15), N0_15_58);
	-- signal N0_15_59 : std_logic;
	PP840 : and2 port map (X(44), Y(15), N0_15_59);
	-- signal N0_15_60 : std_logic;
	PP841 : and2 port map (X(45), Y(15), N0_15_60);
	-- signal N0_15_61 : std_logic;
	PP842 : and2 port map (X(46), Y(15), N0_15_61);
	-- signal N0_15_62 : std_logic;
	PP843 : and2 port map (X(47), Y(15), N0_15_62);
	-- signal N0_15_63 : std_logic;
	PP844 : and2 port map (X(48), Y(15), N0_15_63);
	-- signal N0_15_64 : std_logic;
	PP845 : and2 port map (X(49), Y(15), N0_15_64);
	-- signal N0_15_65 : std_logic;
	PP846 : and2 port map (X(50), Y(15), N0_15_65);
	-- signal N0_15_66 : std_logic;
	PP847 : and2 port map (X(51), Y(15), N0_15_66);
	-- signal N0_15_67 : std_logic;
	PP848 : and2 port map ('1', Y(15), N0_15_67);
	-- signal N0_16_16 : std_logic;
	PP849 : and2 port map (X(0), Y(16), N0_16_16);
	-- signal N0_16_17 : std_logic;
	PP850 : and2 port map (X(1), Y(16), N0_16_17);
	-- signal N0_16_18 : std_logic;
	PP851 : and2 port map (X(2), Y(16), N0_16_18);
	-- signal N0_16_19 : std_logic;
	PP852 : and2 port map (X(3), Y(16), N0_16_19);
	-- signal N0_16_20 : std_logic;
	PP853 : and2 port map (X(4), Y(16), N0_16_20);
	-- signal N0_16_21 : std_logic;
	PP854 : and2 port map (X(5), Y(16), N0_16_21);
	-- signal N0_16_22 : std_logic;
	PP855 : and2 port map (X(6), Y(16), N0_16_22);
	-- signal N0_16_23 : std_logic;
	PP856 : and2 port map (X(7), Y(16), N0_16_23);
	-- signal N0_16_24 : std_logic;
	PP857 : and2 port map (X(8), Y(16), N0_16_24);
	-- signal N0_16_25 : std_logic;
	PP858 : and2 port map (X(9), Y(16), N0_16_25);
	-- signal N0_16_26 : std_logic;
	PP859 : and2 port map (X(10), Y(16), N0_16_26);
	-- signal N0_16_27 : std_logic;
	PP860 : and2 port map (X(11), Y(16), N0_16_27);
	-- signal N0_16_28 : std_logic;
	PP861 : and2 port map (X(12), Y(16), N0_16_28);
	-- signal N0_16_29 : std_logic;
	PP862 : and2 port map (X(13), Y(16), N0_16_29);
	-- signal N0_16_30 : std_logic;
	PP863 : and2 port map (X(14), Y(16), N0_16_30);
	-- signal N0_16_31 : std_logic;
	PP864 : and2 port map (X(15), Y(16), N0_16_31);
	-- signal N0_16_32 : std_logic;
	PP865 : and2 port map (X(16), Y(16), N0_16_32);
	-- signal N0_16_33 : std_logic;
	PP866 : and2 port map (X(17), Y(16), N0_16_33);
	-- signal N0_16_34 : std_logic;
	PP867 : and2 port map (X(18), Y(16), N0_16_34);
	-- signal N0_16_35 : std_logic;
	PP868 : and2 port map (X(19), Y(16), N0_16_35);
	-- signal N0_16_36 : std_logic;
	PP869 : and2 port map (X(20), Y(16), N0_16_36);
	-- signal N0_16_37 : std_logic;
	PP870 : and2 port map (X(21), Y(16), N0_16_37);
	-- signal N0_16_38 : std_logic;
	PP871 : and2 port map (X(22), Y(16), N0_16_38);
	-- signal N0_16_39 : std_logic;
	PP872 : and2 port map (X(23), Y(16), N0_16_39);
	-- signal N0_16_40 : std_logic;
	PP873 : and2 port map (X(24), Y(16), N0_16_40);
	-- signal N0_16_41 : std_logic;
	PP874 : and2 port map (X(25), Y(16), N0_16_41);
	-- signal N0_16_42 : std_logic;
	PP875 : and2 port map (X(26), Y(16), N0_16_42);
	-- signal N0_16_43 : std_logic;
	PP876 : and2 port map (X(27), Y(16), N0_16_43);
	-- signal N0_16_44 : std_logic;
	PP877 : and2 port map (X(28), Y(16), N0_16_44);
	-- signal N0_16_45 : std_logic;
	PP878 : and2 port map (X(29), Y(16), N0_16_45);
	-- signal N0_16_46 : std_logic;
	PP879 : and2 port map (X(30), Y(16), N0_16_46);
	-- signal N0_16_47 : std_logic;
	PP880 : and2 port map (X(31), Y(16), N0_16_47);
	-- signal N0_16_48 : std_logic;
	PP881 : and2 port map (X(32), Y(16), N0_16_48);
	-- signal N0_16_49 : std_logic;
	PP882 : and2 port map (X(33), Y(16), N0_16_49);
	-- signal N0_16_50 : std_logic;
	PP883 : and2 port map (X(34), Y(16), N0_16_50);
	-- signal N0_16_51 : std_logic;
	PP884 : and2 port map (X(35), Y(16), N0_16_51);
	-- signal N0_16_52 : std_logic;
	PP885 : and2 port map (X(36), Y(16), N0_16_52);
	-- signal N0_16_53 : std_logic;
	PP886 : and2 port map (X(37), Y(16), N0_16_53);
	-- signal N0_16_54 : std_logic;
	PP887 : and2 port map (X(38), Y(16), N0_16_54);
	-- signal N0_16_55 : std_logic;
	PP888 : and2 port map (X(39), Y(16), N0_16_55);
	-- signal N0_16_56 : std_logic;
	PP889 : and2 port map (X(40), Y(16), N0_16_56);
	-- signal N0_16_57 : std_logic;
	PP890 : and2 port map (X(41), Y(16), N0_16_57);
	-- signal N0_16_58 : std_logic;
	PP891 : and2 port map (X(42), Y(16), N0_16_58);
	-- signal N0_16_59 : std_logic;
	PP892 : and2 port map (X(43), Y(16), N0_16_59);
	-- signal N0_16_60 : std_logic;
	PP893 : and2 port map (X(44), Y(16), N0_16_60);
	-- signal N0_16_61 : std_logic;
	PP894 : and2 port map (X(45), Y(16), N0_16_61);
	-- signal N0_16_62 : std_logic;
	PP895 : and2 port map (X(46), Y(16), N0_16_62);
	-- signal N0_16_63 : std_logic;
	PP896 : and2 port map (X(47), Y(16), N0_16_63);
	-- signal N0_16_64 : std_logic;
	PP897 : and2 port map (X(48), Y(16), N0_16_64);
	-- signal N0_16_65 : std_logic;
	PP898 : and2 port map (X(49), Y(16), N0_16_65);
	-- signal N0_16_66 : std_logic;
	PP899 : and2 port map (X(50), Y(16), N0_16_66);
	-- signal N0_16_67 : std_logic;
	PP900 : and2 port map (X(51), Y(16), N0_16_67);
	-- signal N0_16_68 : std_logic;
	PP901 : and2 port map ('1', Y(16), N0_16_68);
	-- signal N0_17_17 : std_logic;
	PP902 : and2 port map (X(0), Y(17), N0_17_17);
	-- signal N0_17_18 : std_logic;
	PP903 : and2 port map (X(1), Y(17), N0_17_18);
	-- signal N0_17_19 : std_logic;
	PP904 : and2 port map (X(2), Y(17), N0_17_19);
	-- signal N0_17_20 : std_logic;
	PP905 : and2 port map (X(3), Y(17), N0_17_20);
	-- signal N0_17_21 : std_logic;
	PP906 : and2 port map (X(4), Y(17), N0_17_21);
	-- signal N0_17_22 : std_logic;
	PP907 : and2 port map (X(5), Y(17), N0_17_22);
	-- signal N0_17_23 : std_logic;
	PP908 : and2 port map (X(6), Y(17), N0_17_23);
	-- signal N0_17_24 : std_logic;
	PP909 : and2 port map (X(7), Y(17), N0_17_24);
	-- signal N0_17_25 : std_logic;
	PP910 : and2 port map (X(8), Y(17), N0_17_25);
	-- signal N0_17_26 : std_logic;
	PP911 : and2 port map (X(9), Y(17), N0_17_26);
	-- signal N0_17_27 : std_logic;
	PP912 : and2 port map (X(10), Y(17), N0_17_27);
	-- signal N0_17_28 : std_logic;
	PP913 : and2 port map (X(11), Y(17), N0_17_28);
	-- signal N0_17_29 : std_logic;
	PP914 : and2 port map (X(12), Y(17), N0_17_29);
	-- signal N0_17_30 : std_logic;
	PP915 : and2 port map (X(13), Y(17), N0_17_30);
	-- signal N0_17_31 : std_logic;
	PP916 : and2 port map (X(14), Y(17), N0_17_31);
	-- signal N0_17_32 : std_logic;
	PP917 : and2 port map (X(15), Y(17), N0_17_32);
	-- signal N0_17_33 : std_logic;
	PP918 : and2 port map (X(16), Y(17), N0_17_33);
	-- signal N0_17_34 : std_logic;
	PP919 : and2 port map (X(17), Y(17), N0_17_34);
	-- signal N0_17_35 : std_logic;
	PP920 : and2 port map (X(18), Y(17), N0_17_35);
	-- signal N0_17_36 : std_logic;
	PP921 : and2 port map (X(19), Y(17), N0_17_36);
	-- signal N0_17_37 : std_logic;
	PP922 : and2 port map (X(20), Y(17), N0_17_37);
	-- signal N0_17_38 : std_logic;
	PP923 : and2 port map (X(21), Y(17), N0_17_38);
	-- signal N0_17_39 : std_logic;
	PP924 : and2 port map (X(22), Y(17), N0_17_39);
	-- signal N0_17_40 : std_logic;
	PP925 : and2 port map (X(23), Y(17), N0_17_40);
	-- signal N0_17_41 : std_logic;
	PP926 : and2 port map (X(24), Y(17), N0_17_41);
	-- signal N0_17_42 : std_logic;
	PP927 : and2 port map (X(25), Y(17), N0_17_42);
	-- signal N0_17_43 : std_logic;
	PP928 : and2 port map (X(26), Y(17), N0_17_43);
	-- signal N0_17_44 : std_logic;
	PP929 : and2 port map (X(27), Y(17), N0_17_44);
	-- signal N0_17_45 : std_logic;
	PP930 : and2 port map (X(28), Y(17), N0_17_45);
	-- signal N0_17_46 : std_logic;
	PP931 : and2 port map (X(29), Y(17), N0_17_46);
	-- signal N0_17_47 : std_logic;
	PP932 : and2 port map (X(30), Y(17), N0_17_47);
	-- signal N0_17_48 : std_logic;
	PP933 : and2 port map (X(31), Y(17), N0_17_48);
	-- signal N0_17_49 : std_logic;
	PP934 : and2 port map (X(32), Y(17), N0_17_49);
	-- signal N0_17_50 : std_logic;
	PP935 : and2 port map (X(33), Y(17), N0_17_50);
	-- signal N0_17_51 : std_logic;
	PP936 : and2 port map (X(34), Y(17), N0_17_51);
	-- signal N0_17_52 : std_logic;
	PP937 : and2 port map (X(35), Y(17), N0_17_52);
	-- signal N0_17_53 : std_logic;
	PP938 : and2 port map (X(36), Y(17), N0_17_53);
	-- signal N0_17_54 : std_logic;
	PP939 : and2 port map (X(37), Y(17), N0_17_54);
	-- signal N0_17_55 : std_logic;
	PP940 : and2 port map (X(38), Y(17), N0_17_55);
	-- signal N0_17_56 : std_logic;
	PP941 : and2 port map (X(39), Y(17), N0_17_56);
	-- signal N0_17_57 : std_logic;
	PP942 : and2 port map (X(40), Y(17), N0_17_57);
	-- signal N0_17_58 : std_logic;
	PP943 : and2 port map (X(41), Y(17), N0_17_58);
	-- signal N0_17_59 : std_logic;
	PP944 : and2 port map (X(42), Y(17), N0_17_59);
	-- signal N0_17_60 : std_logic;
	PP945 : and2 port map (X(43), Y(17), N0_17_60);
	-- signal N0_17_61 : std_logic;
	PP946 : and2 port map (X(44), Y(17), N0_17_61);
	-- signal N0_17_62 : std_logic;
	PP947 : and2 port map (X(45), Y(17), N0_17_62);
	-- signal N0_17_63 : std_logic;
	PP948 : and2 port map (X(46), Y(17), N0_17_63);
	-- signal N0_17_64 : std_logic;
	PP949 : and2 port map (X(47), Y(17), N0_17_64);
	-- signal N0_17_65 : std_logic;
	PP950 : and2 port map (X(48), Y(17), N0_17_65);
	-- signal N0_17_66 : std_logic;
	PP951 : and2 port map (X(49), Y(17), N0_17_66);
	-- signal N0_17_67 : std_logic;
	PP952 : and2 port map (X(50), Y(17), N0_17_67);
	-- signal N0_17_68 : std_logic;
	PP953 : and2 port map (X(51), Y(17), N0_17_68);
	-- signal N0_17_69 : std_logic;
	PP954 : and2 port map ('1', Y(17), N0_17_69);
	-- signal N0_18_18 : std_logic;
	PP955 : and2 port map (X(0), Y(18), N0_18_18);
	-- signal N0_18_19 : std_logic;
	PP956 : and2 port map (X(1), Y(18), N0_18_19);
	-- signal N0_18_20 : std_logic;
	PP957 : and2 port map (X(2), Y(18), N0_18_20);
	-- signal N0_18_21 : std_logic;
	PP958 : and2 port map (X(3), Y(18), N0_18_21);
	-- signal N0_18_22 : std_logic;
	PP959 : and2 port map (X(4), Y(18), N0_18_22);
	-- signal N0_18_23 : std_logic;
	PP960 : and2 port map (X(5), Y(18), N0_18_23);
	-- signal N0_18_24 : std_logic;
	PP961 : and2 port map (X(6), Y(18), N0_18_24);
	-- signal N0_18_25 : std_logic;
	PP962 : and2 port map (X(7), Y(18), N0_18_25);
	-- signal N0_18_26 : std_logic;
	PP963 : and2 port map (X(8), Y(18), N0_18_26);
	-- signal N0_18_27 : std_logic;
	PP964 : and2 port map (X(9), Y(18), N0_18_27);
	-- signal N0_18_28 : std_logic;
	PP965 : and2 port map (X(10), Y(18), N0_18_28);
	-- signal N0_18_29 : std_logic;
	PP966 : and2 port map (X(11), Y(18), N0_18_29);
	-- signal N0_18_30 : std_logic;
	PP967 : and2 port map (X(12), Y(18), N0_18_30);
	-- signal N0_18_31 : std_logic;
	PP968 : and2 port map (X(13), Y(18), N0_18_31);
	-- signal N0_18_32 : std_logic;
	PP969 : and2 port map (X(14), Y(18), N0_18_32);
	-- signal N0_18_33 : std_logic;
	PP970 : and2 port map (X(15), Y(18), N0_18_33);
	-- signal N0_18_34 : std_logic;
	PP971 : and2 port map (X(16), Y(18), N0_18_34);
	-- signal N0_18_35 : std_logic;
	PP972 : and2 port map (X(17), Y(18), N0_18_35);
	-- signal N0_18_36 : std_logic;
	PP973 : and2 port map (X(18), Y(18), N0_18_36);
	-- signal N0_18_37 : std_logic;
	PP974 : and2 port map (X(19), Y(18), N0_18_37);
	-- signal N0_18_38 : std_logic;
	PP975 : and2 port map (X(20), Y(18), N0_18_38);
	-- signal N0_18_39 : std_logic;
	PP976 : and2 port map (X(21), Y(18), N0_18_39);
	-- signal N0_18_40 : std_logic;
	PP977 : and2 port map (X(22), Y(18), N0_18_40);
	-- signal N0_18_41 : std_logic;
	PP978 : and2 port map (X(23), Y(18), N0_18_41);
	-- signal N0_18_42 : std_logic;
	PP979 : and2 port map (X(24), Y(18), N0_18_42);
	-- signal N0_18_43 : std_logic;
	PP980 : and2 port map (X(25), Y(18), N0_18_43);
	-- signal N0_18_44 : std_logic;
	PP981 : and2 port map (X(26), Y(18), N0_18_44);
	-- signal N0_18_45 : std_logic;
	PP982 : and2 port map (X(27), Y(18), N0_18_45);
	-- signal N0_18_46 : std_logic;
	PP983 : and2 port map (X(28), Y(18), N0_18_46);
	-- signal N0_18_47 : std_logic;
	PP984 : and2 port map (X(29), Y(18), N0_18_47);
	-- signal N0_18_48 : std_logic;
	PP985 : and2 port map (X(30), Y(18), N0_18_48);
	-- signal N0_18_49 : std_logic;
	PP986 : and2 port map (X(31), Y(18), N0_18_49);
	-- signal N0_18_50 : std_logic;
	PP987 : and2 port map (X(32), Y(18), N0_18_50);
	-- signal N0_18_51 : std_logic;
	PP988 : and2 port map (X(33), Y(18), N0_18_51);
	-- signal N0_18_52 : std_logic;
	PP989 : and2 port map (X(34), Y(18), N0_18_52);
	-- signal N0_18_53 : std_logic;
	PP990 : and2 port map (X(35), Y(18), N0_18_53);
	-- signal N0_18_54 : std_logic;
	PP991 : and2 port map (X(36), Y(18), N0_18_54);
	-- signal N0_18_55 : std_logic;
	PP992 : and2 port map (X(37), Y(18), N0_18_55);
	-- signal N0_18_56 : std_logic;
	PP993 : and2 port map (X(38), Y(18), N0_18_56);
	-- signal N0_18_57 : std_logic;
	PP994 : and2 port map (X(39), Y(18), N0_18_57);
	-- signal N0_18_58 : std_logic;
	PP995 : and2 port map (X(40), Y(18), N0_18_58);
	-- signal N0_18_59 : std_logic;
	PP996 : and2 port map (X(41), Y(18), N0_18_59);
	-- signal N0_18_60 : std_logic;
	PP997 : and2 port map (X(42), Y(18), N0_18_60);
	-- signal N0_18_61 : std_logic;
	PP998 : and2 port map (X(43), Y(18), N0_18_61);
	-- signal N0_18_62 : std_logic;
	PP999 : and2 port map (X(44), Y(18), N0_18_62);
	-- signal N0_18_63 : std_logic;
	PP1000 : and2 port map (X(45), Y(18), N0_18_63);
	-- signal N0_18_64 : std_logic;
	PP1001 : and2 port map (X(46), Y(18), N0_18_64);
	-- signal N0_18_65 : std_logic;
	PP1002 : and2 port map (X(47), Y(18), N0_18_65);
	-- signal N0_18_66 : std_logic;
	PP1003 : and2 port map (X(48), Y(18), N0_18_66);
	-- signal N0_18_67 : std_logic;
	PP1004 : and2 port map (X(49), Y(18), N0_18_67);
	-- signal N0_18_68 : std_logic;
	PP1005 : and2 port map (X(50), Y(18), N0_18_68);
	-- signal N0_18_69 : std_logic;
	PP1006 : and2 port map (X(51), Y(18), N0_18_69);
	-- signal N0_18_70 : std_logic;
	PP1007 : and2 port map ('1', Y(18), N0_18_70);
	-- signal N0_19_19 : std_logic;
	PP1008 : and2 port map (X(0), Y(19), N0_19_19);
	-- signal N0_19_20 : std_logic;
	PP1009 : and2 port map (X(1), Y(19), N0_19_20);
	-- signal N0_19_21 : std_logic;
	PP1010 : and2 port map (X(2), Y(19), N0_19_21);
	-- signal N0_19_22 : std_logic;
	PP1011 : and2 port map (X(3), Y(19), N0_19_22);
	-- signal N0_19_23 : std_logic;
	PP1012 : and2 port map (X(4), Y(19), N0_19_23);
	-- signal N0_19_24 : std_logic;
	PP1013 : and2 port map (X(5), Y(19), N0_19_24);
	-- signal N0_19_25 : std_logic;
	PP1014 : and2 port map (X(6), Y(19), N0_19_25);
	-- signal N0_19_26 : std_logic;
	PP1015 : and2 port map (X(7), Y(19), N0_19_26);
	-- signal N0_19_27 : std_logic;
	PP1016 : and2 port map (X(8), Y(19), N0_19_27);
	-- signal N0_19_28 : std_logic;
	PP1017 : and2 port map (X(9), Y(19), N0_19_28);
	-- signal N0_19_29 : std_logic;
	PP1018 : and2 port map (X(10), Y(19), N0_19_29);
	-- signal N0_19_30 : std_logic;
	PP1019 : and2 port map (X(11), Y(19), N0_19_30);
	-- signal N0_19_31 : std_logic;
	PP1020 : and2 port map (X(12), Y(19), N0_19_31);
	-- signal N0_19_32 : std_logic;
	PP1021 : and2 port map (X(13), Y(19), N0_19_32);
	-- signal N0_19_33 : std_logic;
	PP1022 : and2 port map (X(14), Y(19), N0_19_33);
	-- signal N0_19_34 : std_logic;
	PP1023 : and2 port map (X(15), Y(19), N0_19_34);
	-- signal N0_19_35 : std_logic;
	PP1024 : and2 port map (X(16), Y(19), N0_19_35);
	-- signal N0_19_36 : std_logic;
	PP1025 : and2 port map (X(17), Y(19), N0_19_36);
	-- signal N0_19_37 : std_logic;
	PP1026 : and2 port map (X(18), Y(19), N0_19_37);
	-- signal N0_19_38 : std_logic;
	PP1027 : and2 port map (X(19), Y(19), N0_19_38);
	-- signal N0_19_39 : std_logic;
	PP1028 : and2 port map (X(20), Y(19), N0_19_39);
	-- signal N0_19_40 : std_logic;
	PP1029 : and2 port map (X(21), Y(19), N0_19_40);
	-- signal N0_19_41 : std_logic;
	PP1030 : and2 port map (X(22), Y(19), N0_19_41);
	-- signal N0_19_42 : std_logic;
	PP1031 : and2 port map (X(23), Y(19), N0_19_42);
	-- signal N0_19_43 : std_logic;
	PP1032 : and2 port map (X(24), Y(19), N0_19_43);
	-- signal N0_19_44 : std_logic;
	PP1033 : and2 port map (X(25), Y(19), N0_19_44);
	-- signal N0_19_45 : std_logic;
	PP1034 : and2 port map (X(26), Y(19), N0_19_45);
	-- signal N0_19_46 : std_logic;
	PP1035 : and2 port map (X(27), Y(19), N0_19_46);
	-- signal N0_19_47 : std_logic;
	PP1036 : and2 port map (X(28), Y(19), N0_19_47);
	-- signal N0_19_48 : std_logic;
	PP1037 : and2 port map (X(29), Y(19), N0_19_48);
	-- signal N0_19_49 : std_logic;
	PP1038 : and2 port map (X(30), Y(19), N0_19_49);
	-- signal N0_19_50 : std_logic;
	PP1039 : and2 port map (X(31), Y(19), N0_19_50);
	-- signal N0_19_51 : std_logic;
	PP1040 : and2 port map (X(32), Y(19), N0_19_51);
	-- signal N0_19_52 : std_logic;
	PP1041 : and2 port map (X(33), Y(19), N0_19_52);
	-- signal N0_19_53 : std_logic;
	PP1042 : and2 port map (X(34), Y(19), N0_19_53);
	-- signal N0_19_54 : std_logic;
	PP1043 : and2 port map (X(35), Y(19), N0_19_54);
	-- signal N0_19_55 : std_logic;
	PP1044 : and2 port map (X(36), Y(19), N0_19_55);
	-- signal N0_19_56 : std_logic;
	PP1045 : and2 port map (X(37), Y(19), N0_19_56);
	-- signal N0_19_57 : std_logic;
	PP1046 : and2 port map (X(38), Y(19), N0_19_57);
	-- signal N0_19_58 : std_logic;
	PP1047 : and2 port map (X(39), Y(19), N0_19_58);
	-- signal N0_19_59 : std_logic;
	PP1048 : and2 port map (X(40), Y(19), N0_19_59);
	-- signal N0_19_60 : std_logic;
	PP1049 : and2 port map (X(41), Y(19), N0_19_60);
	-- signal N0_19_61 : std_logic;
	PP1050 : and2 port map (X(42), Y(19), N0_19_61);
	-- signal N0_19_62 : std_logic;
	PP1051 : and2 port map (X(43), Y(19), N0_19_62);
	-- signal N0_19_63 : std_logic;
	PP1052 : and2 port map (X(44), Y(19), N0_19_63);
	-- signal N0_19_64 : std_logic;
	PP1053 : and2 port map (X(45), Y(19), N0_19_64);
	-- signal N0_19_65 : std_logic;
	PP1054 : and2 port map (X(46), Y(19), N0_19_65);
	-- signal N0_19_66 : std_logic;
	PP1055 : and2 port map (X(47), Y(19), N0_19_66);
	-- signal N0_19_67 : std_logic;
	PP1056 : and2 port map (X(48), Y(19), N0_19_67);
	-- signal N0_19_68 : std_logic;
	PP1057 : and2 port map (X(49), Y(19), N0_19_68);
	-- signal N0_19_69 : std_logic;
	PP1058 : and2 port map (X(50), Y(19), N0_19_69);
	-- signal N0_19_70 : std_logic;
	PP1059 : and2 port map (X(51), Y(19), N0_19_70);
	-- signal N0_19_71 : std_logic;
	PP1060 : and2 port map ('1', Y(19), N0_19_71);
	-- signal N0_20_20 : std_logic;
	PP1061 : and2 port map (X(0), Y(20), N0_20_20);
	-- signal N0_20_21 : std_logic;
	PP1062 : and2 port map (X(1), Y(20), N0_20_21);
	-- signal N0_20_22 : std_logic;
	PP1063 : and2 port map (X(2), Y(20), N0_20_22);
	-- signal N0_20_23 : std_logic;
	PP1064 : and2 port map (X(3), Y(20), N0_20_23);
	-- signal N0_20_24 : std_logic;
	PP1065 : and2 port map (X(4), Y(20), N0_20_24);
	-- signal N0_20_25 : std_logic;
	PP1066 : and2 port map (X(5), Y(20), N0_20_25);
	-- signal N0_20_26 : std_logic;
	PP1067 : and2 port map (X(6), Y(20), N0_20_26);
	-- signal N0_20_27 : std_logic;
	PP1068 : and2 port map (X(7), Y(20), N0_20_27);
	-- signal N0_20_28 : std_logic;
	PP1069 : and2 port map (X(8), Y(20), N0_20_28);
	-- signal N0_20_29 : std_logic;
	PP1070 : and2 port map (X(9), Y(20), N0_20_29);
	-- signal N0_20_30 : std_logic;
	PP1071 : and2 port map (X(10), Y(20), N0_20_30);
	-- signal N0_20_31 : std_logic;
	PP1072 : and2 port map (X(11), Y(20), N0_20_31);
	-- signal N0_20_32 : std_logic;
	PP1073 : and2 port map (X(12), Y(20), N0_20_32);
	-- signal N0_20_33 : std_logic;
	PP1074 : and2 port map (X(13), Y(20), N0_20_33);
	-- signal N0_20_34 : std_logic;
	PP1075 : and2 port map (X(14), Y(20), N0_20_34);
	-- signal N0_20_35 : std_logic;
	PP1076 : and2 port map (X(15), Y(20), N0_20_35);
	-- signal N0_20_36 : std_logic;
	PP1077 : and2 port map (X(16), Y(20), N0_20_36);
	-- signal N0_20_37 : std_logic;
	PP1078 : and2 port map (X(17), Y(20), N0_20_37);
	-- signal N0_20_38 : std_logic;
	PP1079 : and2 port map (X(18), Y(20), N0_20_38);
	-- signal N0_20_39 : std_logic;
	PP1080 : and2 port map (X(19), Y(20), N0_20_39);
	-- signal N0_20_40 : std_logic;
	PP1081 : and2 port map (X(20), Y(20), N0_20_40);
	-- signal N0_20_41 : std_logic;
	PP1082 : and2 port map (X(21), Y(20), N0_20_41);
	-- signal N0_20_42 : std_logic;
	PP1083 : and2 port map (X(22), Y(20), N0_20_42);
	-- signal N0_20_43 : std_logic;
	PP1084 : and2 port map (X(23), Y(20), N0_20_43);
	-- signal N0_20_44 : std_logic;
	PP1085 : and2 port map (X(24), Y(20), N0_20_44);
	-- signal N0_20_45 : std_logic;
	PP1086 : and2 port map (X(25), Y(20), N0_20_45);
	-- signal N0_20_46 : std_logic;
	PP1087 : and2 port map (X(26), Y(20), N0_20_46);
	-- signal N0_20_47 : std_logic;
	PP1088 : and2 port map (X(27), Y(20), N0_20_47);
	-- signal N0_20_48 : std_logic;
	PP1089 : and2 port map (X(28), Y(20), N0_20_48);
	-- signal N0_20_49 : std_logic;
	PP1090 : and2 port map (X(29), Y(20), N0_20_49);
	-- signal N0_20_50 : std_logic;
	PP1091 : and2 port map (X(30), Y(20), N0_20_50);
	-- signal N0_20_51 : std_logic;
	PP1092 : and2 port map (X(31), Y(20), N0_20_51);
	-- signal N0_20_52 : std_logic;
	PP1093 : and2 port map (X(32), Y(20), N0_20_52);
	-- signal N0_20_53 : std_logic;
	PP1094 : and2 port map (X(33), Y(20), N0_20_53);
	-- signal N0_20_54 : std_logic;
	PP1095 : and2 port map (X(34), Y(20), N0_20_54);
	-- signal N0_20_55 : std_logic;
	PP1096 : and2 port map (X(35), Y(20), N0_20_55);
	-- signal N0_20_56 : std_logic;
	PP1097 : and2 port map (X(36), Y(20), N0_20_56);
	-- signal N0_20_57 : std_logic;
	PP1098 : and2 port map (X(37), Y(20), N0_20_57);
	-- signal N0_20_58 : std_logic;
	PP1099 : and2 port map (X(38), Y(20), N0_20_58);
	-- signal N0_20_59 : std_logic;
	PP1100 : and2 port map (X(39), Y(20), N0_20_59);
	-- signal N0_20_60 : std_logic;
	PP1101 : and2 port map (X(40), Y(20), N0_20_60);
	-- signal N0_20_61 : std_logic;
	PP1102 : and2 port map (X(41), Y(20), N0_20_61);
	-- signal N0_20_62 : std_logic;
	PP1103 : and2 port map (X(42), Y(20), N0_20_62);
	-- signal N0_20_63 : std_logic;
	PP1104 : and2 port map (X(43), Y(20), N0_20_63);
	-- signal N0_20_64 : std_logic;
	PP1105 : and2 port map (X(44), Y(20), N0_20_64);
	-- signal N0_20_65 : std_logic;
	PP1106 : and2 port map (X(45), Y(20), N0_20_65);
	-- signal N0_20_66 : std_logic;
	PP1107 : and2 port map (X(46), Y(20), N0_20_66);
	-- signal N0_20_67 : std_logic;
	PP1108 : and2 port map (X(47), Y(20), N0_20_67);
	-- signal N0_20_68 : std_logic;
	PP1109 : and2 port map (X(48), Y(20), N0_20_68);
	-- signal N0_20_69 : std_logic;
	PP1110 : and2 port map (X(49), Y(20), N0_20_69);
	-- signal N0_20_70 : std_logic;
	PP1111 : and2 port map (X(50), Y(20), N0_20_70);
	-- signal N0_20_71 : std_logic;
	PP1112 : and2 port map (X(51), Y(20), N0_20_71);
	-- signal N0_20_72 : std_logic;
	PP1113 : and2 port map ('1', Y(20), N0_20_72);
	-- signal N0_21_21 : std_logic;
	PP1114 : and2 port map (X(0), Y(21), N0_21_21);
	-- signal N0_21_22 : std_logic;
	PP1115 : and2 port map (X(1), Y(21), N0_21_22);
	-- signal N0_21_23 : std_logic;
	PP1116 : and2 port map (X(2), Y(21), N0_21_23);
	-- signal N0_21_24 : std_logic;
	PP1117 : and2 port map (X(3), Y(21), N0_21_24);
	-- signal N0_21_25 : std_logic;
	PP1118 : and2 port map (X(4), Y(21), N0_21_25);
	-- signal N0_21_26 : std_logic;
	PP1119 : and2 port map (X(5), Y(21), N0_21_26);
	-- signal N0_21_27 : std_logic;
	PP1120 : and2 port map (X(6), Y(21), N0_21_27);
	-- signal N0_21_28 : std_logic;
	PP1121 : and2 port map (X(7), Y(21), N0_21_28);
	-- signal N0_21_29 : std_logic;
	PP1122 : and2 port map (X(8), Y(21), N0_21_29);
	-- signal N0_21_30 : std_logic;
	PP1123 : and2 port map (X(9), Y(21), N0_21_30);
	-- signal N0_21_31 : std_logic;
	PP1124 : and2 port map (X(10), Y(21), N0_21_31);
	-- signal N0_21_32 : std_logic;
	PP1125 : and2 port map (X(11), Y(21), N0_21_32);
	-- signal N0_21_33 : std_logic;
	PP1126 : and2 port map (X(12), Y(21), N0_21_33);
	-- signal N0_21_34 : std_logic;
	PP1127 : and2 port map (X(13), Y(21), N0_21_34);
	-- signal N0_21_35 : std_logic;
	PP1128 : and2 port map (X(14), Y(21), N0_21_35);
	-- signal N0_21_36 : std_logic;
	PP1129 : and2 port map (X(15), Y(21), N0_21_36);
	-- signal N0_21_37 : std_logic;
	PP1130 : and2 port map (X(16), Y(21), N0_21_37);
	-- signal N0_21_38 : std_logic;
	PP1131 : and2 port map (X(17), Y(21), N0_21_38);
	-- signal N0_21_39 : std_logic;
	PP1132 : and2 port map (X(18), Y(21), N0_21_39);
	-- signal N0_21_40 : std_logic;
	PP1133 : and2 port map (X(19), Y(21), N0_21_40);
	-- signal N0_21_41 : std_logic;
	PP1134 : and2 port map (X(20), Y(21), N0_21_41);
	-- signal N0_21_42 : std_logic;
	PP1135 : and2 port map (X(21), Y(21), N0_21_42);
	-- signal N0_21_43 : std_logic;
	PP1136 : and2 port map (X(22), Y(21), N0_21_43);
	-- signal N0_21_44 : std_logic;
	PP1137 : and2 port map (X(23), Y(21), N0_21_44);
	-- signal N0_21_45 : std_logic;
	PP1138 : and2 port map (X(24), Y(21), N0_21_45);
	-- signal N0_21_46 : std_logic;
	PP1139 : and2 port map (X(25), Y(21), N0_21_46);
	-- signal N0_21_47 : std_logic;
	PP1140 : and2 port map (X(26), Y(21), N0_21_47);
	-- signal N0_21_48 : std_logic;
	PP1141 : and2 port map (X(27), Y(21), N0_21_48);
	-- signal N0_21_49 : std_logic;
	PP1142 : and2 port map (X(28), Y(21), N0_21_49);
	-- signal N0_21_50 : std_logic;
	PP1143 : and2 port map (X(29), Y(21), N0_21_50);
	-- signal N0_21_51 : std_logic;
	PP1144 : and2 port map (X(30), Y(21), N0_21_51);
	-- signal N0_21_52 : std_logic;
	PP1145 : and2 port map (X(31), Y(21), N0_21_52);
	-- signal N0_21_53 : std_logic;
	PP1146 : and2 port map (X(32), Y(21), N0_21_53);
	-- signal N0_21_54 : std_logic;
	PP1147 : and2 port map (X(33), Y(21), N0_21_54);
	-- signal N0_21_55 : std_logic;
	PP1148 : and2 port map (X(34), Y(21), N0_21_55);
	-- signal N0_21_56 : std_logic;
	PP1149 : and2 port map (X(35), Y(21), N0_21_56);
	-- signal N0_21_57 : std_logic;
	PP1150 : and2 port map (X(36), Y(21), N0_21_57);
	-- signal N0_21_58 : std_logic;
	PP1151 : and2 port map (X(37), Y(21), N0_21_58);
	-- signal N0_21_59 : std_logic;
	PP1152 : and2 port map (X(38), Y(21), N0_21_59);
	-- signal N0_21_60 : std_logic;
	PP1153 : and2 port map (X(39), Y(21), N0_21_60);
	-- signal N0_21_61 : std_logic;
	PP1154 : and2 port map (X(40), Y(21), N0_21_61);
	-- signal N0_21_62 : std_logic;
	PP1155 : and2 port map (X(41), Y(21), N0_21_62);
	-- signal N0_21_63 : std_logic;
	PP1156 : and2 port map (X(42), Y(21), N0_21_63);
	-- signal N0_21_64 : std_logic;
	PP1157 : and2 port map (X(43), Y(21), N0_21_64);
	-- signal N0_21_65 : std_logic;
	PP1158 : and2 port map (X(44), Y(21), N0_21_65);
	-- signal N0_21_66 : std_logic;
	PP1159 : and2 port map (X(45), Y(21), N0_21_66);
	-- signal N0_21_67 : std_logic;
	PP1160 : and2 port map (X(46), Y(21), N0_21_67);
	-- signal N0_21_68 : std_logic;
	PP1161 : and2 port map (X(47), Y(21), N0_21_68);
	-- signal N0_21_69 : std_logic;
	PP1162 : and2 port map (X(48), Y(21), N0_21_69);
	-- signal N0_21_70 : std_logic;
	PP1163 : and2 port map (X(49), Y(21), N0_21_70);
	-- signal N0_21_71 : std_logic;
	PP1164 : and2 port map (X(50), Y(21), N0_21_71);
	-- signal N0_21_72 : std_logic;
	PP1165 : and2 port map (X(51), Y(21), N0_21_72);
	-- signal N0_21_73 : std_logic;
	PP1166 : and2 port map ('1', Y(21), N0_21_73);
	-- signal N0_22_22 : std_logic;
	PP1167 : and2 port map (X(0), Y(22), N0_22_22);
	-- signal N0_22_23 : std_logic;
	PP1168 : and2 port map (X(1), Y(22), N0_22_23);
	-- signal N0_22_24 : std_logic;
	PP1169 : and2 port map (X(2), Y(22), N0_22_24);
	-- signal N0_22_25 : std_logic;
	PP1170 : and2 port map (X(3), Y(22), N0_22_25);
	-- signal N0_22_26 : std_logic;
	PP1171 : and2 port map (X(4), Y(22), N0_22_26);
	-- signal N0_22_27 : std_logic;
	PP1172 : and2 port map (X(5), Y(22), N0_22_27);
	-- signal N0_22_28 : std_logic;
	PP1173 : and2 port map (X(6), Y(22), N0_22_28);
	-- signal N0_22_29 : std_logic;
	PP1174 : and2 port map (X(7), Y(22), N0_22_29);
	-- signal N0_22_30 : std_logic;
	PP1175 : and2 port map (X(8), Y(22), N0_22_30);
	-- signal N0_22_31 : std_logic;
	PP1176 : and2 port map (X(9), Y(22), N0_22_31);
	-- signal N0_22_32 : std_logic;
	PP1177 : and2 port map (X(10), Y(22), N0_22_32);
	-- signal N0_22_33 : std_logic;
	PP1178 : and2 port map (X(11), Y(22), N0_22_33);
	-- signal N0_22_34 : std_logic;
	PP1179 : and2 port map (X(12), Y(22), N0_22_34);
	-- signal N0_22_35 : std_logic;
	PP1180 : and2 port map (X(13), Y(22), N0_22_35);
	-- signal N0_22_36 : std_logic;
	PP1181 : and2 port map (X(14), Y(22), N0_22_36);
	-- signal N0_22_37 : std_logic;
	PP1182 : and2 port map (X(15), Y(22), N0_22_37);
	-- signal N0_22_38 : std_logic;
	PP1183 : and2 port map (X(16), Y(22), N0_22_38);
	-- signal N0_22_39 : std_logic;
	PP1184 : and2 port map (X(17), Y(22), N0_22_39);
	-- signal N0_22_40 : std_logic;
	PP1185 : and2 port map (X(18), Y(22), N0_22_40);
	-- signal N0_22_41 : std_logic;
	PP1186 : and2 port map (X(19), Y(22), N0_22_41);
	-- signal N0_22_42 : std_logic;
	PP1187 : and2 port map (X(20), Y(22), N0_22_42);
	-- signal N0_22_43 : std_logic;
	PP1188 : and2 port map (X(21), Y(22), N0_22_43);
	-- signal N0_22_44 : std_logic;
	PP1189 : and2 port map (X(22), Y(22), N0_22_44);
	-- signal N0_22_45 : std_logic;
	PP1190 : and2 port map (X(23), Y(22), N0_22_45);
	-- signal N0_22_46 : std_logic;
	PP1191 : and2 port map (X(24), Y(22), N0_22_46);
	-- signal N0_22_47 : std_logic;
	PP1192 : and2 port map (X(25), Y(22), N0_22_47);
	-- signal N0_22_48 : std_logic;
	PP1193 : and2 port map (X(26), Y(22), N0_22_48);
	-- signal N0_22_49 : std_logic;
	PP1194 : and2 port map (X(27), Y(22), N0_22_49);
	-- signal N0_22_50 : std_logic;
	PP1195 : and2 port map (X(28), Y(22), N0_22_50);
	-- signal N0_22_51 : std_logic;
	PP1196 : and2 port map (X(29), Y(22), N0_22_51);
	-- signal N0_22_52 : std_logic;
	PP1197 : and2 port map (X(30), Y(22), N0_22_52);
	-- signal N0_22_53 : std_logic;
	PP1198 : and2 port map (X(31), Y(22), N0_22_53);
	-- signal N0_22_54 : std_logic;
	PP1199 : and2 port map (X(32), Y(22), N0_22_54);
	-- signal N0_22_55 : std_logic;
	PP1200 : and2 port map (X(33), Y(22), N0_22_55);
	-- signal N0_22_56 : std_logic;
	PP1201 : and2 port map (X(34), Y(22), N0_22_56);
	-- signal N0_22_57 : std_logic;
	PP1202 : and2 port map (X(35), Y(22), N0_22_57);
	-- signal N0_22_58 : std_logic;
	PP1203 : and2 port map (X(36), Y(22), N0_22_58);
	-- signal N0_22_59 : std_logic;
	PP1204 : and2 port map (X(37), Y(22), N0_22_59);
	-- signal N0_22_60 : std_logic;
	PP1205 : and2 port map (X(38), Y(22), N0_22_60);
	-- signal N0_22_61 : std_logic;
	PP1206 : and2 port map (X(39), Y(22), N0_22_61);
	-- signal N0_22_62 : std_logic;
	PP1207 : and2 port map (X(40), Y(22), N0_22_62);
	-- signal N0_22_63 : std_logic;
	PP1208 : and2 port map (X(41), Y(22), N0_22_63);
	-- signal N0_22_64 : std_logic;
	PP1209 : and2 port map (X(42), Y(22), N0_22_64);
	-- signal N0_22_65 : std_logic;
	PP1210 : and2 port map (X(43), Y(22), N0_22_65);
	-- signal N0_22_66 : std_logic;
	PP1211 : and2 port map (X(44), Y(22), N0_22_66);
	-- signal N0_22_67 : std_logic;
	PP1212 : and2 port map (X(45), Y(22), N0_22_67);
	-- signal N0_22_68 : std_logic;
	PP1213 : and2 port map (X(46), Y(22), N0_22_68);
	-- signal N0_22_69 : std_logic;
	PP1214 : and2 port map (X(47), Y(22), N0_22_69);
	-- signal N0_22_70 : std_logic;
	PP1215 : and2 port map (X(48), Y(22), N0_22_70);
	-- signal N0_22_71 : std_logic;
	PP1216 : and2 port map (X(49), Y(22), N0_22_71);
	-- signal N0_22_72 : std_logic;
	PP1217 : and2 port map (X(50), Y(22), N0_22_72);
	-- signal N0_22_73 : std_logic;
	PP1218 : and2 port map (X(51), Y(22), N0_22_73);
	-- signal N0_22_74 : std_logic;
	PP1219 : and2 port map ('1', Y(22), N0_22_74);
	-- signal N0_23_23 : std_logic;
	PP1220 : and2 port map (X(0), Y(23), N0_23_23);
	-- signal N0_23_24 : std_logic;
	PP1221 : and2 port map (X(1), Y(23), N0_23_24);
	-- signal N0_23_25 : std_logic;
	PP1222 : and2 port map (X(2), Y(23), N0_23_25);
	-- signal N0_23_26 : std_logic;
	PP1223 : and2 port map (X(3), Y(23), N0_23_26);
	-- signal N0_23_27 : std_logic;
	PP1224 : and2 port map (X(4), Y(23), N0_23_27);
	-- signal N0_23_28 : std_logic;
	PP1225 : and2 port map (X(5), Y(23), N0_23_28);
	-- signal N0_23_29 : std_logic;
	PP1226 : and2 port map (X(6), Y(23), N0_23_29);
	-- signal N0_23_30 : std_logic;
	PP1227 : and2 port map (X(7), Y(23), N0_23_30);
	-- signal N0_23_31 : std_logic;
	PP1228 : and2 port map (X(8), Y(23), N0_23_31);
	-- signal N0_23_32 : std_logic;
	PP1229 : and2 port map (X(9), Y(23), N0_23_32);
	-- signal N0_23_33 : std_logic;
	PP1230 : and2 port map (X(10), Y(23), N0_23_33);
	-- signal N0_23_34 : std_logic;
	PP1231 : and2 port map (X(11), Y(23), N0_23_34);
	-- signal N0_23_35 : std_logic;
	PP1232 : and2 port map (X(12), Y(23), N0_23_35);
	-- signal N0_23_36 : std_logic;
	PP1233 : and2 port map (X(13), Y(23), N0_23_36);
	-- signal N0_23_37 : std_logic;
	PP1234 : and2 port map (X(14), Y(23), N0_23_37);
	-- signal N0_23_38 : std_logic;
	PP1235 : and2 port map (X(15), Y(23), N0_23_38);
	-- signal N0_23_39 : std_logic;
	PP1236 : and2 port map (X(16), Y(23), N0_23_39);
	-- signal N0_23_40 : std_logic;
	PP1237 : and2 port map (X(17), Y(23), N0_23_40);
	-- signal N0_23_41 : std_logic;
	PP1238 : and2 port map (X(18), Y(23), N0_23_41);
	-- signal N0_23_42 : std_logic;
	PP1239 : and2 port map (X(19), Y(23), N0_23_42);
	-- signal N0_23_43 : std_logic;
	PP1240 : and2 port map (X(20), Y(23), N0_23_43);
	-- signal N0_23_44 : std_logic;
	PP1241 : and2 port map (X(21), Y(23), N0_23_44);
	-- signal N0_23_45 : std_logic;
	PP1242 : and2 port map (X(22), Y(23), N0_23_45);
	-- signal N0_23_46 : std_logic;
	PP1243 : and2 port map (X(23), Y(23), N0_23_46);
	-- signal N0_23_47 : std_logic;
	PP1244 : and2 port map (X(24), Y(23), N0_23_47);
	-- signal N0_23_48 : std_logic;
	PP1245 : and2 port map (X(25), Y(23), N0_23_48);
	-- signal N0_23_49 : std_logic;
	PP1246 : and2 port map (X(26), Y(23), N0_23_49);
	-- signal N0_23_50 : std_logic;
	PP1247 : and2 port map (X(27), Y(23), N0_23_50);
	-- signal N0_23_51 : std_logic;
	PP1248 : and2 port map (X(28), Y(23), N0_23_51);
	-- signal N0_23_52 : std_logic;
	PP1249 : and2 port map (X(29), Y(23), N0_23_52);
	-- signal N0_23_53 : std_logic;
	PP1250 : and2 port map (X(30), Y(23), N0_23_53);
	-- signal N0_23_54 : std_logic;
	PP1251 : and2 port map (X(31), Y(23), N0_23_54);
	-- signal N0_23_55 : std_logic;
	PP1252 : and2 port map (X(32), Y(23), N0_23_55);
	-- signal N0_23_56 : std_logic;
	PP1253 : and2 port map (X(33), Y(23), N0_23_56);
	-- signal N0_23_57 : std_logic;
	PP1254 : and2 port map (X(34), Y(23), N0_23_57);
	-- signal N0_23_58 : std_logic;
	PP1255 : and2 port map (X(35), Y(23), N0_23_58);
	-- signal N0_23_59 : std_logic;
	PP1256 : and2 port map (X(36), Y(23), N0_23_59);
	-- signal N0_23_60 : std_logic;
	PP1257 : and2 port map (X(37), Y(23), N0_23_60);
	-- signal N0_23_61 : std_logic;
	PP1258 : and2 port map (X(38), Y(23), N0_23_61);
	-- signal N0_23_62 : std_logic;
	PP1259 : and2 port map (X(39), Y(23), N0_23_62);
	-- signal N0_23_63 : std_logic;
	PP1260 : and2 port map (X(40), Y(23), N0_23_63);
	-- signal N0_23_64 : std_logic;
	PP1261 : and2 port map (X(41), Y(23), N0_23_64);
	-- signal N0_23_65 : std_logic;
	PP1262 : and2 port map (X(42), Y(23), N0_23_65);
	-- signal N0_23_66 : std_logic;
	PP1263 : and2 port map (X(43), Y(23), N0_23_66);
	-- signal N0_23_67 : std_logic;
	PP1264 : and2 port map (X(44), Y(23), N0_23_67);
	-- signal N0_23_68 : std_logic;
	PP1265 : and2 port map (X(45), Y(23), N0_23_68);
	-- signal N0_23_69 : std_logic;
	PP1266 : and2 port map (X(46), Y(23), N0_23_69);
	-- signal N0_23_70 : std_logic;
	PP1267 : and2 port map (X(47), Y(23), N0_23_70);
	-- signal N0_23_71 : std_logic;
	PP1268 : and2 port map (X(48), Y(23), N0_23_71);
	-- signal N0_23_72 : std_logic;
	PP1269 : and2 port map (X(49), Y(23), N0_23_72);
	-- signal N0_23_73 : std_logic;
	PP1270 : and2 port map (X(50), Y(23), N0_23_73);
	-- signal N0_23_74 : std_logic;
	PP1271 : and2 port map (X(51), Y(23), N0_23_74);
	-- signal N0_23_75 : std_logic;
	PP1272 : and2 port map ('1', Y(23), N0_23_75);
	-- signal N0_24_24 : std_logic;
	PP1273 : and2 port map (X(0), Y(24), N0_24_24);
	-- signal N0_24_25 : std_logic;
	PP1274 : and2 port map (X(1), Y(24), N0_24_25);
	-- signal N0_24_26 : std_logic;
	PP1275 : and2 port map (X(2), Y(24), N0_24_26);
	-- signal N0_24_27 : std_logic;
	PP1276 : and2 port map (X(3), Y(24), N0_24_27);
	-- signal N0_24_28 : std_logic;
	PP1277 : and2 port map (X(4), Y(24), N0_24_28);
	-- signal N0_24_29 : std_logic;
	PP1278 : and2 port map (X(5), Y(24), N0_24_29);
	-- signal N0_24_30 : std_logic;
	PP1279 : and2 port map (X(6), Y(24), N0_24_30);
	-- signal N0_24_31 : std_logic;
	PP1280 : and2 port map (X(7), Y(24), N0_24_31);
	-- signal N0_24_32 : std_logic;
	PP1281 : and2 port map (X(8), Y(24), N0_24_32);
	-- signal N0_24_33 : std_logic;
	PP1282 : and2 port map (X(9), Y(24), N0_24_33);
	-- signal N0_24_34 : std_logic;
	PP1283 : and2 port map (X(10), Y(24), N0_24_34);
	-- signal N0_24_35 : std_logic;
	PP1284 : and2 port map (X(11), Y(24), N0_24_35);
	-- signal N0_24_36 : std_logic;
	PP1285 : and2 port map (X(12), Y(24), N0_24_36);
	-- signal N0_24_37 : std_logic;
	PP1286 : and2 port map (X(13), Y(24), N0_24_37);
	-- signal N0_24_38 : std_logic;
	PP1287 : and2 port map (X(14), Y(24), N0_24_38);
	-- signal N0_24_39 : std_logic;
	PP1288 : and2 port map (X(15), Y(24), N0_24_39);
	-- signal N0_24_40 : std_logic;
	PP1289 : and2 port map (X(16), Y(24), N0_24_40);
	-- signal N0_24_41 : std_logic;
	PP1290 : and2 port map (X(17), Y(24), N0_24_41);
	-- signal N0_24_42 : std_logic;
	PP1291 : and2 port map (X(18), Y(24), N0_24_42);
	-- signal N0_24_43 : std_logic;
	PP1292 : and2 port map (X(19), Y(24), N0_24_43);
	-- signal N0_24_44 : std_logic;
	PP1293 : and2 port map (X(20), Y(24), N0_24_44);
	-- signal N0_24_45 : std_logic;
	PP1294 : and2 port map (X(21), Y(24), N0_24_45);
	-- signal N0_24_46 : std_logic;
	PP1295 : and2 port map (X(22), Y(24), N0_24_46);
	-- signal N0_24_47 : std_logic;
	PP1296 : and2 port map (X(23), Y(24), N0_24_47);
	-- signal N0_24_48 : std_logic;
	PP1297 : and2 port map (X(24), Y(24), N0_24_48);
	-- signal N0_24_49 : std_logic;
	PP1298 : and2 port map (X(25), Y(24), N0_24_49);
	-- signal N0_24_50 : std_logic;
	PP1299 : and2 port map (X(26), Y(24), N0_24_50);
	-- signal N0_24_51 : std_logic;
	PP1300 : and2 port map (X(27), Y(24), N0_24_51);
	-- signal N0_24_52 : std_logic;
	PP1301 : and2 port map (X(28), Y(24), N0_24_52);
	-- signal N0_24_53 : std_logic;
	PP1302 : and2 port map (X(29), Y(24), N0_24_53);
	-- signal N0_24_54 : std_logic;
	PP1303 : and2 port map (X(30), Y(24), N0_24_54);
	-- signal N0_24_55 : std_logic;
	PP1304 : and2 port map (X(31), Y(24), N0_24_55);
	-- signal N0_24_56 : std_logic;
	PP1305 : and2 port map (X(32), Y(24), N0_24_56);
	-- signal N0_24_57 : std_logic;
	PP1306 : and2 port map (X(33), Y(24), N0_24_57);
	-- signal N0_24_58 : std_logic;
	PP1307 : and2 port map (X(34), Y(24), N0_24_58);
	-- signal N0_24_59 : std_logic;
	PP1308 : and2 port map (X(35), Y(24), N0_24_59);
	-- signal N0_24_60 : std_logic;
	PP1309 : and2 port map (X(36), Y(24), N0_24_60);
	-- signal N0_24_61 : std_logic;
	PP1310 : and2 port map (X(37), Y(24), N0_24_61);
	-- signal N0_24_62 : std_logic;
	PP1311 : and2 port map (X(38), Y(24), N0_24_62);
	-- signal N0_24_63 : std_logic;
	PP1312 : and2 port map (X(39), Y(24), N0_24_63);
	-- signal N0_24_64 : std_logic;
	PP1313 : and2 port map (X(40), Y(24), N0_24_64);
	-- signal N0_24_65 : std_logic;
	PP1314 : and2 port map (X(41), Y(24), N0_24_65);
	-- signal N0_24_66 : std_logic;
	PP1315 : and2 port map (X(42), Y(24), N0_24_66);
	-- signal N0_24_67 : std_logic;
	PP1316 : and2 port map (X(43), Y(24), N0_24_67);
	-- signal N0_24_68 : std_logic;
	PP1317 : and2 port map (X(44), Y(24), N0_24_68);
	-- signal N0_24_69 : std_logic;
	PP1318 : and2 port map (X(45), Y(24), N0_24_69);
	-- signal N0_24_70 : std_logic;
	PP1319 : and2 port map (X(46), Y(24), N0_24_70);
	-- signal N0_24_71 : std_logic;
	PP1320 : and2 port map (X(47), Y(24), N0_24_71);
	-- signal N0_24_72 : std_logic;
	PP1321 : and2 port map (X(48), Y(24), N0_24_72);
	-- signal N0_24_73 : std_logic;
	PP1322 : and2 port map (X(49), Y(24), N0_24_73);
	-- signal N0_24_74 : std_logic;
	PP1323 : and2 port map (X(50), Y(24), N0_24_74);
	-- signal N0_24_75 : std_logic;
	PP1324 : and2 port map (X(51), Y(24), N0_24_75);
	-- signal N0_24_76 : std_logic;
	PP1325 : and2 port map ('1', Y(24), N0_24_76);
	-- signal N0_25_25 : std_logic;
	PP1326 : and2 port map (X(0), Y(25), N0_25_25);
	-- signal N0_25_26 : std_logic;
	PP1327 : and2 port map (X(1), Y(25), N0_25_26);
	-- signal N0_25_27 : std_logic;
	PP1328 : and2 port map (X(2), Y(25), N0_25_27);
	-- signal N0_25_28 : std_logic;
	PP1329 : and2 port map (X(3), Y(25), N0_25_28);
	-- signal N0_25_29 : std_logic;
	PP1330 : and2 port map (X(4), Y(25), N0_25_29);
	-- signal N0_25_30 : std_logic;
	PP1331 : and2 port map (X(5), Y(25), N0_25_30);
	-- signal N0_25_31 : std_logic;
	PP1332 : and2 port map (X(6), Y(25), N0_25_31);
	-- signal N0_25_32 : std_logic;
	PP1333 : and2 port map (X(7), Y(25), N0_25_32);
	-- signal N0_25_33 : std_logic;
	PP1334 : and2 port map (X(8), Y(25), N0_25_33);
	-- signal N0_25_34 : std_logic;
	PP1335 : and2 port map (X(9), Y(25), N0_25_34);
	-- signal N0_25_35 : std_logic;
	PP1336 : and2 port map (X(10), Y(25), N0_25_35);
	-- signal N0_25_36 : std_logic;
	PP1337 : and2 port map (X(11), Y(25), N0_25_36);
	-- signal N0_25_37 : std_logic;
	PP1338 : and2 port map (X(12), Y(25), N0_25_37);
	-- signal N0_25_38 : std_logic;
	PP1339 : and2 port map (X(13), Y(25), N0_25_38);
	-- signal N0_25_39 : std_logic;
	PP1340 : and2 port map (X(14), Y(25), N0_25_39);
	-- signal N0_25_40 : std_logic;
	PP1341 : and2 port map (X(15), Y(25), N0_25_40);
	-- signal N0_25_41 : std_logic;
	PP1342 : and2 port map (X(16), Y(25), N0_25_41);
	-- signal N0_25_42 : std_logic;
	PP1343 : and2 port map (X(17), Y(25), N0_25_42);
	-- signal N0_25_43 : std_logic;
	PP1344 : and2 port map (X(18), Y(25), N0_25_43);
	-- signal N0_25_44 : std_logic;
	PP1345 : and2 port map (X(19), Y(25), N0_25_44);
	-- signal N0_25_45 : std_logic;
	PP1346 : and2 port map (X(20), Y(25), N0_25_45);
	-- signal N0_25_46 : std_logic;
	PP1347 : and2 port map (X(21), Y(25), N0_25_46);
	-- signal N0_25_47 : std_logic;
	PP1348 : and2 port map (X(22), Y(25), N0_25_47);
	-- signal N0_25_48 : std_logic;
	PP1349 : and2 port map (X(23), Y(25), N0_25_48);
	-- signal N0_25_49 : std_logic;
	PP1350 : and2 port map (X(24), Y(25), N0_25_49);
	-- signal N0_25_50 : std_logic;
	PP1351 : and2 port map (X(25), Y(25), N0_25_50);
	-- signal N0_25_51 : std_logic;
	PP1352 : and2 port map (X(26), Y(25), N0_25_51);
	-- signal N0_25_52 : std_logic;
	PP1353 : and2 port map (X(27), Y(25), N0_25_52);
	-- signal N0_25_53 : std_logic;
	PP1354 : and2 port map (X(28), Y(25), N0_25_53);
	-- signal N0_25_54 : std_logic;
	PP1355 : and2 port map (X(29), Y(25), N0_25_54);
	-- signal N0_25_55 : std_logic;
	PP1356 : and2 port map (X(30), Y(25), N0_25_55);
	-- signal N0_25_56 : std_logic;
	PP1357 : and2 port map (X(31), Y(25), N0_25_56);
	-- signal N0_25_57 : std_logic;
	PP1358 : and2 port map (X(32), Y(25), N0_25_57);
	-- signal N0_25_58 : std_logic;
	PP1359 : and2 port map (X(33), Y(25), N0_25_58);
	-- signal N0_25_59 : std_logic;
	PP1360 : and2 port map (X(34), Y(25), N0_25_59);
	-- signal N0_25_60 : std_logic;
	PP1361 : and2 port map (X(35), Y(25), N0_25_60);
	-- signal N0_25_61 : std_logic;
	PP1362 : and2 port map (X(36), Y(25), N0_25_61);
	-- signal N0_25_62 : std_logic;
	PP1363 : and2 port map (X(37), Y(25), N0_25_62);
	-- signal N0_25_63 : std_logic;
	PP1364 : and2 port map (X(38), Y(25), N0_25_63);
	-- signal N0_25_64 : std_logic;
	PP1365 : and2 port map (X(39), Y(25), N0_25_64);
	-- signal N0_25_65 : std_logic;
	PP1366 : and2 port map (X(40), Y(25), N0_25_65);
	-- signal N0_25_66 : std_logic;
	PP1367 : and2 port map (X(41), Y(25), N0_25_66);
	-- signal N0_25_67 : std_logic;
	PP1368 : and2 port map (X(42), Y(25), N0_25_67);
	-- signal N0_25_68 : std_logic;
	PP1369 : and2 port map (X(43), Y(25), N0_25_68);
	-- signal N0_25_69 : std_logic;
	PP1370 : and2 port map (X(44), Y(25), N0_25_69);
	-- signal N0_25_70 : std_logic;
	PP1371 : and2 port map (X(45), Y(25), N0_25_70);
	-- signal N0_25_71 : std_logic;
	PP1372 : and2 port map (X(46), Y(25), N0_25_71);
	-- signal N0_25_72 : std_logic;
	PP1373 : and2 port map (X(47), Y(25), N0_25_72);
	-- signal N0_25_73 : std_logic;
	PP1374 : and2 port map (X(48), Y(25), N0_25_73);
	-- signal N0_25_74 : std_logic;
	PP1375 : and2 port map (X(49), Y(25), N0_25_74);
	-- signal N0_25_75 : std_logic;
	PP1376 : and2 port map (X(50), Y(25), N0_25_75);
	-- signal N0_25_76 : std_logic;
	PP1377 : and2 port map (X(51), Y(25), N0_25_76);
	-- signal N0_25_77 : std_logic;
	PP1378 : and2 port map ('1', Y(25), N0_25_77);
	-- signal N0_26_26 : std_logic;
	PP1379 : and2 port map (X(0), Y(26), N0_26_26);
	-- signal N0_26_27 : std_logic;
	PP1380 : and2 port map (X(1), Y(26), N0_26_27);
	-- signal N0_26_28 : std_logic;
	PP1381 : and2 port map (X(2), Y(26), N0_26_28);
	-- signal N0_26_29 : std_logic;
	PP1382 : and2 port map (X(3), Y(26), N0_26_29);
	-- signal N0_26_30 : std_logic;
	PP1383 : and2 port map (X(4), Y(26), N0_26_30);
	-- signal N0_26_31 : std_logic;
	PP1384 : and2 port map (X(5), Y(26), N0_26_31);
	-- signal N0_26_32 : std_logic;
	PP1385 : and2 port map (X(6), Y(26), N0_26_32);
	-- signal N0_26_33 : std_logic;
	PP1386 : and2 port map (X(7), Y(26), N0_26_33);
	-- signal N0_26_34 : std_logic;
	PP1387 : and2 port map (X(8), Y(26), N0_26_34);
	-- signal N0_26_35 : std_logic;
	PP1388 : and2 port map (X(9), Y(26), N0_26_35);
	-- signal N0_26_36 : std_logic;
	PP1389 : and2 port map (X(10), Y(26), N0_26_36);
	-- signal N0_26_37 : std_logic;
	PP1390 : and2 port map (X(11), Y(26), N0_26_37);
	-- signal N0_26_38 : std_logic;
	PP1391 : and2 port map (X(12), Y(26), N0_26_38);
	-- signal N0_26_39 : std_logic;
	PP1392 : and2 port map (X(13), Y(26), N0_26_39);
	-- signal N0_26_40 : std_logic;
	PP1393 : and2 port map (X(14), Y(26), N0_26_40);
	-- signal N0_26_41 : std_logic;
	PP1394 : and2 port map (X(15), Y(26), N0_26_41);
	-- signal N0_26_42 : std_logic;
	PP1395 : and2 port map (X(16), Y(26), N0_26_42);
	-- signal N0_26_43 : std_logic;
	PP1396 : and2 port map (X(17), Y(26), N0_26_43);
	-- signal N0_26_44 : std_logic;
	PP1397 : and2 port map (X(18), Y(26), N0_26_44);
	-- signal N0_26_45 : std_logic;
	PP1398 : and2 port map (X(19), Y(26), N0_26_45);
	-- signal N0_26_46 : std_logic;
	PP1399 : and2 port map (X(20), Y(26), N0_26_46);
	-- signal N0_26_47 : std_logic;
	PP1400 : and2 port map (X(21), Y(26), N0_26_47);
	-- signal N0_26_48 : std_logic;
	PP1401 : and2 port map (X(22), Y(26), N0_26_48);
	-- signal N0_26_49 : std_logic;
	PP1402 : and2 port map (X(23), Y(26), N0_26_49);
	-- signal N0_26_50 : std_logic;
	PP1403 : and2 port map (X(24), Y(26), N0_26_50);
	-- signal N0_26_51 : std_logic;
	PP1404 : and2 port map (X(25), Y(26), N0_26_51);
	-- signal N0_26_52 : std_logic;
	PP1405 : and2 port map (X(26), Y(26), N0_26_52);
	-- signal N0_26_53 : std_logic;
	PP1406 : and2 port map (X(27), Y(26), N0_26_53);
	-- signal N0_26_54 : std_logic;
	PP1407 : and2 port map (X(28), Y(26), N0_26_54);
	-- signal N0_26_55 : std_logic;
	PP1408 : and2 port map (X(29), Y(26), N0_26_55);
	-- signal N0_26_56 : std_logic;
	PP1409 : and2 port map (X(30), Y(26), N0_26_56);
	-- signal N0_26_57 : std_logic;
	PP1410 : and2 port map (X(31), Y(26), N0_26_57);
	-- signal N0_26_58 : std_logic;
	PP1411 : and2 port map (X(32), Y(26), N0_26_58);
	-- signal N0_26_59 : std_logic;
	PP1412 : and2 port map (X(33), Y(26), N0_26_59);
	-- signal N0_26_60 : std_logic;
	PP1413 : and2 port map (X(34), Y(26), N0_26_60);
	-- signal N0_26_61 : std_logic;
	PP1414 : and2 port map (X(35), Y(26), N0_26_61);
	-- signal N0_26_62 : std_logic;
	PP1415 : and2 port map (X(36), Y(26), N0_26_62);
	-- signal N0_26_63 : std_logic;
	PP1416 : and2 port map (X(37), Y(26), N0_26_63);
	-- signal N0_26_64 : std_logic;
	PP1417 : and2 port map (X(38), Y(26), N0_26_64);
	-- signal N0_26_65 : std_logic;
	PP1418 : and2 port map (X(39), Y(26), N0_26_65);
	-- signal N0_26_66 : std_logic;
	PP1419 : and2 port map (X(40), Y(26), N0_26_66);
	-- signal N0_26_67 : std_logic;
	PP1420 : and2 port map (X(41), Y(26), N0_26_67);
	-- signal N0_26_68 : std_logic;
	PP1421 : and2 port map (X(42), Y(26), N0_26_68);
	-- signal N0_26_69 : std_logic;
	PP1422 : and2 port map (X(43), Y(26), N0_26_69);
	-- signal N0_26_70 : std_logic;
	PP1423 : and2 port map (X(44), Y(26), N0_26_70);
	-- signal N0_26_71 : std_logic;
	PP1424 : and2 port map (X(45), Y(26), N0_26_71);
	-- signal N0_26_72 : std_logic;
	PP1425 : and2 port map (X(46), Y(26), N0_26_72);
	-- signal N0_26_73 : std_logic;
	PP1426 : and2 port map (X(47), Y(26), N0_26_73);
	-- signal N0_26_74 : std_logic;
	PP1427 : and2 port map (X(48), Y(26), N0_26_74);
	-- signal N0_26_75 : std_logic;
	PP1428 : and2 port map (X(49), Y(26), N0_26_75);
	-- signal N0_26_76 : std_logic;
	PP1429 : and2 port map (X(50), Y(26), N0_26_76);
	-- signal N0_26_77 : std_logic;
	PP1430 : and2 port map (X(51), Y(26), N0_26_77);
	-- signal N0_26_78 : std_logic;
	PP1431 : and2 port map ('1', Y(26), N0_26_78);
	-- signal N0_27_27 : std_logic;
	PP1432 : and2 port map (X(0), Y(27), N0_27_27);
	-- signal N0_27_28 : std_logic;
	PP1433 : and2 port map (X(1), Y(27), N0_27_28);
	-- signal N0_27_29 : std_logic;
	PP1434 : and2 port map (X(2), Y(27), N0_27_29);
	-- signal N0_27_30 : std_logic;
	PP1435 : and2 port map (X(3), Y(27), N0_27_30);
	-- signal N0_27_31 : std_logic;
	PP1436 : and2 port map (X(4), Y(27), N0_27_31);
	-- signal N0_27_32 : std_logic;
	PP1437 : and2 port map (X(5), Y(27), N0_27_32);
	-- signal N0_27_33 : std_logic;
	PP1438 : and2 port map (X(6), Y(27), N0_27_33);
	-- signal N0_27_34 : std_logic;
	PP1439 : and2 port map (X(7), Y(27), N0_27_34);
	-- signal N0_27_35 : std_logic;
	PP1440 : and2 port map (X(8), Y(27), N0_27_35);
	-- signal N0_27_36 : std_logic;
	PP1441 : and2 port map (X(9), Y(27), N0_27_36);
	-- signal N0_27_37 : std_logic;
	PP1442 : and2 port map (X(10), Y(27), N0_27_37);
	-- signal N0_27_38 : std_logic;
	PP1443 : and2 port map (X(11), Y(27), N0_27_38);
	-- signal N0_27_39 : std_logic;
	PP1444 : and2 port map (X(12), Y(27), N0_27_39);
	-- signal N0_27_40 : std_logic;
	PP1445 : and2 port map (X(13), Y(27), N0_27_40);
	-- signal N0_27_41 : std_logic;
	PP1446 : and2 port map (X(14), Y(27), N0_27_41);
	-- signal N0_27_42 : std_logic;
	PP1447 : and2 port map (X(15), Y(27), N0_27_42);
	-- signal N0_27_43 : std_logic;
	PP1448 : and2 port map (X(16), Y(27), N0_27_43);
	-- signal N0_27_44 : std_logic;
	PP1449 : and2 port map (X(17), Y(27), N0_27_44);
	-- signal N0_27_45 : std_logic;
	PP1450 : and2 port map (X(18), Y(27), N0_27_45);
	-- signal N0_27_46 : std_logic;
	PP1451 : and2 port map (X(19), Y(27), N0_27_46);
	-- signal N0_27_47 : std_logic;
	PP1452 : and2 port map (X(20), Y(27), N0_27_47);
	-- signal N0_27_48 : std_logic;
	PP1453 : and2 port map (X(21), Y(27), N0_27_48);
	-- signal N0_27_49 : std_logic;
	PP1454 : and2 port map (X(22), Y(27), N0_27_49);
	-- signal N0_27_50 : std_logic;
	PP1455 : and2 port map (X(23), Y(27), N0_27_50);
	-- signal N0_27_51 : std_logic;
	PP1456 : and2 port map (X(24), Y(27), N0_27_51);
	-- signal N0_27_52 : std_logic;
	PP1457 : and2 port map (X(25), Y(27), N0_27_52);
	-- signal N0_27_53 : std_logic;
	PP1458 : and2 port map (X(26), Y(27), N0_27_53);
	-- signal N0_27_54 : std_logic;
	PP1459 : and2 port map (X(27), Y(27), N0_27_54);
	-- signal N0_27_55 : std_logic;
	PP1460 : and2 port map (X(28), Y(27), N0_27_55);
	-- signal N0_27_56 : std_logic;
	PP1461 : and2 port map (X(29), Y(27), N0_27_56);
	-- signal N0_27_57 : std_logic;
	PP1462 : and2 port map (X(30), Y(27), N0_27_57);
	-- signal N0_27_58 : std_logic;
	PP1463 : and2 port map (X(31), Y(27), N0_27_58);
	-- signal N0_27_59 : std_logic;
	PP1464 : and2 port map (X(32), Y(27), N0_27_59);
	-- signal N0_27_60 : std_logic;
	PP1465 : and2 port map (X(33), Y(27), N0_27_60);
	-- signal N0_27_61 : std_logic;
	PP1466 : and2 port map (X(34), Y(27), N0_27_61);
	-- signal N0_27_62 : std_logic;
	PP1467 : and2 port map (X(35), Y(27), N0_27_62);
	-- signal N0_27_63 : std_logic;
	PP1468 : and2 port map (X(36), Y(27), N0_27_63);
	-- signal N0_27_64 : std_logic;
	PP1469 : and2 port map (X(37), Y(27), N0_27_64);
	-- signal N0_27_65 : std_logic;
	PP1470 : and2 port map (X(38), Y(27), N0_27_65);
	-- signal N0_27_66 : std_logic;
	PP1471 : and2 port map (X(39), Y(27), N0_27_66);
	-- signal N0_27_67 : std_logic;
	PP1472 : and2 port map (X(40), Y(27), N0_27_67);
	-- signal N0_27_68 : std_logic;
	PP1473 : and2 port map (X(41), Y(27), N0_27_68);
	-- signal N0_27_69 : std_logic;
	PP1474 : and2 port map (X(42), Y(27), N0_27_69);
	-- signal N0_27_70 : std_logic;
	PP1475 : and2 port map (X(43), Y(27), N0_27_70);
	-- signal N0_27_71 : std_logic;
	PP1476 : and2 port map (X(44), Y(27), N0_27_71);
	-- signal N0_27_72 : std_logic;
	PP1477 : and2 port map (X(45), Y(27), N0_27_72);
	-- signal N0_27_73 : std_logic;
	PP1478 : and2 port map (X(46), Y(27), N0_27_73);
	-- signal N0_27_74 : std_logic;
	PP1479 : and2 port map (X(47), Y(27), N0_27_74);
	-- signal N0_27_75 : std_logic;
	PP1480 : and2 port map (X(48), Y(27), N0_27_75);
	-- signal N0_27_76 : std_logic;
	PP1481 : and2 port map (X(49), Y(27), N0_27_76);
	-- signal N0_27_77 : std_logic;
	PP1482 : and2 port map (X(50), Y(27), N0_27_77);
	-- signal N0_27_78 : std_logic;
	PP1483 : and2 port map (X(51), Y(27), N0_27_78);
	-- signal N0_27_79 : std_logic;
	PP1484 : and2 port map ('1', Y(27), N0_27_79);
	-- signal N0_28_28 : std_logic;
	PP1485 : and2 port map (X(0), Y(28), N0_28_28);
	-- signal N0_28_29 : std_logic;
	PP1486 : and2 port map (X(1), Y(28), N0_28_29);
	-- signal N0_28_30 : std_logic;
	PP1487 : and2 port map (X(2), Y(28), N0_28_30);
	-- signal N0_28_31 : std_logic;
	PP1488 : and2 port map (X(3), Y(28), N0_28_31);
	-- signal N0_28_32 : std_logic;
	PP1489 : and2 port map (X(4), Y(28), N0_28_32);
	-- signal N0_28_33 : std_logic;
	PP1490 : and2 port map (X(5), Y(28), N0_28_33);
	-- signal N0_28_34 : std_logic;
	PP1491 : and2 port map (X(6), Y(28), N0_28_34);
	-- signal N0_28_35 : std_logic;
	PP1492 : and2 port map (X(7), Y(28), N0_28_35);
	-- signal N0_28_36 : std_logic;
	PP1493 : and2 port map (X(8), Y(28), N0_28_36);
	-- signal N0_28_37 : std_logic;
	PP1494 : and2 port map (X(9), Y(28), N0_28_37);
	-- signal N0_28_38 : std_logic;
	PP1495 : and2 port map (X(10), Y(28), N0_28_38);
	-- signal N0_28_39 : std_logic;
	PP1496 : and2 port map (X(11), Y(28), N0_28_39);
	-- signal N0_28_40 : std_logic;
	PP1497 : and2 port map (X(12), Y(28), N0_28_40);
	-- signal N0_28_41 : std_logic;
	PP1498 : and2 port map (X(13), Y(28), N0_28_41);
	-- signal N0_28_42 : std_logic;
	PP1499 : and2 port map (X(14), Y(28), N0_28_42);
	-- signal N0_28_43 : std_logic;
	PP1500 : and2 port map (X(15), Y(28), N0_28_43);
	-- signal N0_28_44 : std_logic;
	PP1501 : and2 port map (X(16), Y(28), N0_28_44);
	-- signal N0_28_45 : std_logic;
	PP1502 : and2 port map (X(17), Y(28), N0_28_45);
	-- signal N0_28_46 : std_logic;
	PP1503 : and2 port map (X(18), Y(28), N0_28_46);
	-- signal N0_28_47 : std_logic;
	PP1504 : and2 port map (X(19), Y(28), N0_28_47);
	-- signal N0_28_48 : std_logic;
	PP1505 : and2 port map (X(20), Y(28), N0_28_48);
	-- signal N0_28_49 : std_logic;
	PP1506 : and2 port map (X(21), Y(28), N0_28_49);
	-- signal N0_28_50 : std_logic;
	PP1507 : and2 port map (X(22), Y(28), N0_28_50);
	-- signal N0_28_51 : std_logic;
	PP1508 : and2 port map (X(23), Y(28), N0_28_51);
	-- signal N0_28_52 : std_logic;
	PP1509 : and2 port map (X(24), Y(28), N0_28_52);
	-- signal N0_28_53 : std_logic;
	PP1510 : and2 port map (X(25), Y(28), N0_28_53);
	-- signal N0_28_54 : std_logic;
	PP1511 : and2 port map (X(26), Y(28), N0_28_54);
	-- signal N0_28_55 : std_logic;
	PP1512 : and2 port map (X(27), Y(28), N0_28_55);
	-- signal N0_28_56 : std_logic;
	PP1513 : and2 port map (X(28), Y(28), N0_28_56);
	-- signal N0_28_57 : std_logic;
	PP1514 : and2 port map (X(29), Y(28), N0_28_57);
	-- signal N0_28_58 : std_logic;
	PP1515 : and2 port map (X(30), Y(28), N0_28_58);
	-- signal N0_28_59 : std_logic;
	PP1516 : and2 port map (X(31), Y(28), N0_28_59);
	-- signal N0_28_60 : std_logic;
	PP1517 : and2 port map (X(32), Y(28), N0_28_60);
	-- signal N0_28_61 : std_logic;
	PP1518 : and2 port map (X(33), Y(28), N0_28_61);
	-- signal N0_28_62 : std_logic;
	PP1519 : and2 port map (X(34), Y(28), N0_28_62);
	-- signal N0_28_63 : std_logic;
	PP1520 : and2 port map (X(35), Y(28), N0_28_63);
	-- signal N0_28_64 : std_logic;
	PP1521 : and2 port map (X(36), Y(28), N0_28_64);
	-- signal N0_28_65 : std_logic;
	PP1522 : and2 port map (X(37), Y(28), N0_28_65);
	-- signal N0_28_66 : std_logic;
	PP1523 : and2 port map (X(38), Y(28), N0_28_66);
	-- signal N0_28_67 : std_logic;
	PP1524 : and2 port map (X(39), Y(28), N0_28_67);
	-- signal N0_28_68 : std_logic;
	PP1525 : and2 port map (X(40), Y(28), N0_28_68);
	-- signal N0_28_69 : std_logic;
	PP1526 : and2 port map (X(41), Y(28), N0_28_69);
	-- signal N0_28_70 : std_logic;
	PP1527 : and2 port map (X(42), Y(28), N0_28_70);
	-- signal N0_28_71 : std_logic;
	PP1528 : and2 port map (X(43), Y(28), N0_28_71);
	-- signal N0_28_72 : std_logic;
	PP1529 : and2 port map (X(44), Y(28), N0_28_72);
	-- signal N0_28_73 : std_logic;
	PP1530 : and2 port map (X(45), Y(28), N0_28_73);
	-- signal N0_28_74 : std_logic;
	PP1531 : and2 port map (X(46), Y(28), N0_28_74);
	-- signal N0_28_75 : std_logic;
	PP1532 : and2 port map (X(47), Y(28), N0_28_75);
	-- signal N0_28_76 : std_logic;
	PP1533 : and2 port map (X(48), Y(28), N0_28_76);
	-- signal N0_28_77 : std_logic;
	PP1534 : and2 port map (X(49), Y(28), N0_28_77);
	-- signal N0_28_78 : std_logic;
	PP1535 : and2 port map (X(50), Y(28), N0_28_78);
	-- signal N0_28_79 : std_logic;
	PP1536 : and2 port map (X(51), Y(28), N0_28_79);
	-- signal N0_28_80 : std_logic;
	PP1537 : and2 port map ('1', Y(28), N0_28_80);
	-- signal N0_29_29 : std_logic;
	PP1538 : and2 port map (X(0), Y(29), N0_29_29);
	-- signal N0_29_30 : std_logic;
	PP1539 : and2 port map (X(1), Y(29), N0_29_30);
	-- signal N0_29_31 : std_logic;
	PP1540 : and2 port map (X(2), Y(29), N0_29_31);
	-- signal N0_29_32 : std_logic;
	PP1541 : and2 port map (X(3), Y(29), N0_29_32);
	-- signal N0_29_33 : std_logic;
	PP1542 : and2 port map (X(4), Y(29), N0_29_33);
	-- signal N0_29_34 : std_logic;
	PP1543 : and2 port map (X(5), Y(29), N0_29_34);
	-- signal N0_29_35 : std_logic;
	PP1544 : and2 port map (X(6), Y(29), N0_29_35);
	-- signal N0_29_36 : std_logic;
	PP1545 : and2 port map (X(7), Y(29), N0_29_36);
	-- signal N0_29_37 : std_logic;
	PP1546 : and2 port map (X(8), Y(29), N0_29_37);
	-- signal N0_29_38 : std_logic;
	PP1547 : and2 port map (X(9), Y(29), N0_29_38);
	-- signal N0_29_39 : std_logic;
	PP1548 : and2 port map (X(10), Y(29), N0_29_39);
	-- signal N0_29_40 : std_logic;
	PP1549 : and2 port map (X(11), Y(29), N0_29_40);
	-- signal N0_29_41 : std_logic;
	PP1550 : and2 port map (X(12), Y(29), N0_29_41);
	-- signal N0_29_42 : std_logic;
	PP1551 : and2 port map (X(13), Y(29), N0_29_42);
	-- signal N0_29_43 : std_logic;
	PP1552 : and2 port map (X(14), Y(29), N0_29_43);
	-- signal N0_29_44 : std_logic;
	PP1553 : and2 port map (X(15), Y(29), N0_29_44);
	-- signal N0_29_45 : std_logic;
	PP1554 : and2 port map (X(16), Y(29), N0_29_45);
	-- signal N0_29_46 : std_logic;
	PP1555 : and2 port map (X(17), Y(29), N0_29_46);
	-- signal N0_29_47 : std_logic;
	PP1556 : and2 port map (X(18), Y(29), N0_29_47);
	-- signal N0_29_48 : std_logic;
	PP1557 : and2 port map (X(19), Y(29), N0_29_48);
	-- signal N0_29_49 : std_logic;
	PP1558 : and2 port map (X(20), Y(29), N0_29_49);
	-- signal N0_29_50 : std_logic;
	PP1559 : and2 port map (X(21), Y(29), N0_29_50);
	-- signal N0_29_51 : std_logic;
	PP1560 : and2 port map (X(22), Y(29), N0_29_51);
	-- signal N0_29_52 : std_logic;
	PP1561 : and2 port map (X(23), Y(29), N0_29_52);
	-- signal N0_29_53 : std_logic;
	PP1562 : and2 port map (X(24), Y(29), N0_29_53);
	-- signal N0_29_54 : std_logic;
	PP1563 : and2 port map (X(25), Y(29), N0_29_54);
	-- signal N0_29_55 : std_logic;
	PP1564 : and2 port map (X(26), Y(29), N0_29_55);
	-- signal N0_29_56 : std_logic;
	PP1565 : and2 port map (X(27), Y(29), N0_29_56);
	-- signal N0_29_57 : std_logic;
	PP1566 : and2 port map (X(28), Y(29), N0_29_57);
	-- signal N0_29_58 : std_logic;
	PP1567 : and2 port map (X(29), Y(29), N0_29_58);
	-- signal N0_29_59 : std_logic;
	PP1568 : and2 port map (X(30), Y(29), N0_29_59);
	-- signal N0_29_60 : std_logic;
	PP1569 : and2 port map (X(31), Y(29), N0_29_60);
	-- signal N0_29_61 : std_logic;
	PP1570 : and2 port map (X(32), Y(29), N0_29_61);
	-- signal N0_29_62 : std_logic;
	PP1571 : and2 port map (X(33), Y(29), N0_29_62);
	-- signal N0_29_63 : std_logic;
	PP1572 : and2 port map (X(34), Y(29), N0_29_63);
	-- signal N0_29_64 : std_logic;
	PP1573 : and2 port map (X(35), Y(29), N0_29_64);
	-- signal N0_29_65 : std_logic;
	PP1574 : and2 port map (X(36), Y(29), N0_29_65);
	-- signal N0_29_66 : std_logic;
	PP1575 : and2 port map (X(37), Y(29), N0_29_66);
	-- signal N0_29_67 : std_logic;
	PP1576 : and2 port map (X(38), Y(29), N0_29_67);
	-- signal N0_29_68 : std_logic;
	PP1577 : and2 port map (X(39), Y(29), N0_29_68);
	-- signal N0_29_69 : std_logic;
	PP1578 : and2 port map (X(40), Y(29), N0_29_69);
	-- signal N0_29_70 : std_logic;
	PP1579 : and2 port map (X(41), Y(29), N0_29_70);
	-- signal N0_29_71 : std_logic;
	PP1580 : and2 port map (X(42), Y(29), N0_29_71);
	-- signal N0_29_72 : std_logic;
	PP1581 : and2 port map (X(43), Y(29), N0_29_72);
	-- signal N0_29_73 : std_logic;
	PP1582 : and2 port map (X(44), Y(29), N0_29_73);
	-- signal N0_29_74 : std_logic;
	PP1583 : and2 port map (X(45), Y(29), N0_29_74);
	-- signal N0_29_75 : std_logic;
	PP1584 : and2 port map (X(46), Y(29), N0_29_75);
	-- signal N0_29_76 : std_logic;
	PP1585 : and2 port map (X(47), Y(29), N0_29_76);
	-- signal N0_29_77 : std_logic;
	PP1586 : and2 port map (X(48), Y(29), N0_29_77);
	-- signal N0_29_78 : std_logic;
	PP1587 : and2 port map (X(49), Y(29), N0_29_78);
	-- signal N0_29_79 : std_logic;
	PP1588 : and2 port map (X(50), Y(29), N0_29_79);
	-- signal N0_29_80 : std_logic;
	PP1589 : and2 port map (X(51), Y(29), N0_29_80);
	-- signal N0_29_81 : std_logic;
	PP1590 : and2 port map ('1', Y(29), N0_29_81);
	-- signal N0_30_30 : std_logic;
	PP1591 : and2 port map (X(0), Y(30), N0_30_30);
	-- signal N0_30_31 : std_logic;
	PP1592 : and2 port map (X(1), Y(30), N0_30_31);
	-- signal N0_30_32 : std_logic;
	PP1593 : and2 port map (X(2), Y(30), N0_30_32);
	-- signal N0_30_33 : std_logic;
	PP1594 : and2 port map (X(3), Y(30), N0_30_33);
	-- signal N0_30_34 : std_logic;
	PP1595 : and2 port map (X(4), Y(30), N0_30_34);
	-- signal N0_30_35 : std_logic;
	PP1596 : and2 port map (X(5), Y(30), N0_30_35);
	-- signal N0_30_36 : std_logic;
	PP1597 : and2 port map (X(6), Y(30), N0_30_36);
	-- signal N0_30_37 : std_logic;
	PP1598 : and2 port map (X(7), Y(30), N0_30_37);
	-- signal N0_30_38 : std_logic;
	PP1599 : and2 port map (X(8), Y(30), N0_30_38);
	-- signal N0_30_39 : std_logic;
	PP1600 : and2 port map (X(9), Y(30), N0_30_39);
	-- signal N0_30_40 : std_logic;
	PP1601 : and2 port map (X(10), Y(30), N0_30_40);
	-- signal N0_30_41 : std_logic;
	PP1602 : and2 port map (X(11), Y(30), N0_30_41);
	-- signal N0_30_42 : std_logic;
	PP1603 : and2 port map (X(12), Y(30), N0_30_42);
	-- signal N0_30_43 : std_logic;
	PP1604 : and2 port map (X(13), Y(30), N0_30_43);
	-- signal N0_30_44 : std_logic;
	PP1605 : and2 port map (X(14), Y(30), N0_30_44);
	-- signal N0_30_45 : std_logic;
	PP1606 : and2 port map (X(15), Y(30), N0_30_45);
	-- signal N0_30_46 : std_logic;
	PP1607 : and2 port map (X(16), Y(30), N0_30_46);
	-- signal N0_30_47 : std_logic;
	PP1608 : and2 port map (X(17), Y(30), N0_30_47);
	-- signal N0_30_48 : std_logic;
	PP1609 : and2 port map (X(18), Y(30), N0_30_48);
	-- signal N0_30_49 : std_logic;
	PP1610 : and2 port map (X(19), Y(30), N0_30_49);
	-- signal N0_30_50 : std_logic;
	PP1611 : and2 port map (X(20), Y(30), N0_30_50);
	-- signal N0_30_51 : std_logic;
	PP1612 : and2 port map (X(21), Y(30), N0_30_51);
	-- signal N0_30_52 : std_logic;
	PP1613 : and2 port map (X(22), Y(30), N0_30_52);
	-- signal N0_30_53 : std_logic;
	PP1614 : and2 port map (X(23), Y(30), N0_30_53);
	-- signal N0_30_54 : std_logic;
	PP1615 : and2 port map (X(24), Y(30), N0_30_54);
	-- signal N0_30_55 : std_logic;
	PP1616 : and2 port map (X(25), Y(30), N0_30_55);
	-- signal N0_30_56 : std_logic;
	PP1617 : and2 port map (X(26), Y(30), N0_30_56);
	-- signal N0_30_57 : std_logic;
	PP1618 : and2 port map (X(27), Y(30), N0_30_57);
	-- signal N0_30_58 : std_logic;
	PP1619 : and2 port map (X(28), Y(30), N0_30_58);
	-- signal N0_30_59 : std_logic;
	PP1620 : and2 port map (X(29), Y(30), N0_30_59);
	-- signal N0_30_60 : std_logic;
	PP1621 : and2 port map (X(30), Y(30), N0_30_60);
	-- signal N0_30_61 : std_logic;
	PP1622 : and2 port map (X(31), Y(30), N0_30_61);
	-- signal N0_30_62 : std_logic;
	PP1623 : and2 port map (X(32), Y(30), N0_30_62);
	-- signal N0_30_63 : std_logic;
	PP1624 : and2 port map (X(33), Y(30), N0_30_63);
	-- signal N0_30_64 : std_logic;
	PP1625 : and2 port map (X(34), Y(30), N0_30_64);
	-- signal N0_30_65 : std_logic;
	PP1626 : and2 port map (X(35), Y(30), N0_30_65);
	-- signal N0_30_66 : std_logic;
	PP1627 : and2 port map (X(36), Y(30), N0_30_66);
	-- signal N0_30_67 : std_logic;
	PP1628 : and2 port map (X(37), Y(30), N0_30_67);
	-- signal N0_30_68 : std_logic;
	PP1629 : and2 port map (X(38), Y(30), N0_30_68);
	-- signal N0_30_69 : std_logic;
	PP1630 : and2 port map (X(39), Y(30), N0_30_69);
	-- signal N0_30_70 : std_logic;
	PP1631 : and2 port map (X(40), Y(30), N0_30_70);
	-- signal N0_30_71 : std_logic;
	PP1632 : and2 port map (X(41), Y(30), N0_30_71);
	-- signal N0_30_72 : std_logic;
	PP1633 : and2 port map (X(42), Y(30), N0_30_72);
	-- signal N0_30_73 : std_logic;
	PP1634 : and2 port map (X(43), Y(30), N0_30_73);
	-- signal N0_30_74 : std_logic;
	PP1635 : and2 port map (X(44), Y(30), N0_30_74);
	-- signal N0_30_75 : std_logic;
	PP1636 : and2 port map (X(45), Y(30), N0_30_75);
	-- signal N0_30_76 : std_logic;
	PP1637 : and2 port map (X(46), Y(30), N0_30_76);
	-- signal N0_30_77 : std_logic;
	PP1638 : and2 port map (X(47), Y(30), N0_30_77);
	-- signal N0_30_78 : std_logic;
	PP1639 : and2 port map (X(48), Y(30), N0_30_78);
	-- signal N0_30_79 : std_logic;
	PP1640 : and2 port map (X(49), Y(30), N0_30_79);
	-- signal N0_30_80 : std_logic;
	PP1641 : and2 port map (X(50), Y(30), N0_30_80);
	-- signal N0_30_81 : std_logic;
	PP1642 : and2 port map (X(51), Y(30), N0_30_81);
	-- signal N0_30_82 : std_logic;
	PP1643 : and2 port map ('1', Y(30), N0_30_82);
	-- signal N0_31_31 : std_logic;
	PP1644 : and2 port map (X(0), Y(31), N0_31_31);
	-- signal N0_31_32 : std_logic;
	PP1645 : and2 port map (X(1), Y(31), N0_31_32);
	-- signal N0_31_33 : std_logic;
	PP1646 : and2 port map (X(2), Y(31), N0_31_33);
	-- signal N0_31_34 : std_logic;
	PP1647 : and2 port map (X(3), Y(31), N0_31_34);
	-- signal N0_31_35 : std_logic;
	PP1648 : and2 port map (X(4), Y(31), N0_31_35);
	-- signal N0_31_36 : std_logic;
	PP1649 : and2 port map (X(5), Y(31), N0_31_36);
	-- signal N0_31_37 : std_logic;
	PP1650 : and2 port map (X(6), Y(31), N0_31_37);
	-- signal N0_31_38 : std_logic;
	PP1651 : and2 port map (X(7), Y(31), N0_31_38);
	-- signal N0_31_39 : std_logic;
	PP1652 : and2 port map (X(8), Y(31), N0_31_39);
	-- signal N0_31_40 : std_logic;
	PP1653 : and2 port map (X(9), Y(31), N0_31_40);
	-- signal N0_31_41 : std_logic;
	PP1654 : and2 port map (X(10), Y(31), N0_31_41);
	-- signal N0_31_42 : std_logic;
	PP1655 : and2 port map (X(11), Y(31), N0_31_42);
	-- signal N0_31_43 : std_logic;
	PP1656 : and2 port map (X(12), Y(31), N0_31_43);
	-- signal N0_31_44 : std_logic;
	PP1657 : and2 port map (X(13), Y(31), N0_31_44);
	-- signal N0_31_45 : std_logic;
	PP1658 : and2 port map (X(14), Y(31), N0_31_45);
	-- signal N0_31_46 : std_logic;
	PP1659 : and2 port map (X(15), Y(31), N0_31_46);
	-- signal N0_31_47 : std_logic;
	PP1660 : and2 port map (X(16), Y(31), N0_31_47);
	-- signal N0_31_48 : std_logic;
	PP1661 : and2 port map (X(17), Y(31), N0_31_48);
	-- signal N0_31_49 : std_logic;
	PP1662 : and2 port map (X(18), Y(31), N0_31_49);
	-- signal N0_31_50 : std_logic;
	PP1663 : and2 port map (X(19), Y(31), N0_31_50);
	-- signal N0_31_51 : std_logic;
	PP1664 : and2 port map (X(20), Y(31), N0_31_51);
	-- signal N0_31_52 : std_logic;
	PP1665 : and2 port map (X(21), Y(31), N0_31_52);
	-- signal N0_31_53 : std_logic;
	PP1666 : and2 port map (X(22), Y(31), N0_31_53);
	-- signal N0_31_54 : std_logic;
	PP1667 : and2 port map (X(23), Y(31), N0_31_54);
	-- signal N0_31_55 : std_logic;
	PP1668 : and2 port map (X(24), Y(31), N0_31_55);
	-- signal N0_31_56 : std_logic;
	PP1669 : and2 port map (X(25), Y(31), N0_31_56);
	-- signal N0_31_57 : std_logic;
	PP1670 : and2 port map (X(26), Y(31), N0_31_57);
	-- signal N0_31_58 : std_logic;
	PP1671 : and2 port map (X(27), Y(31), N0_31_58);
	-- signal N0_31_59 : std_logic;
	PP1672 : and2 port map (X(28), Y(31), N0_31_59);
	-- signal N0_31_60 : std_logic;
	PP1673 : and2 port map (X(29), Y(31), N0_31_60);
	-- signal N0_31_61 : std_logic;
	PP1674 : and2 port map (X(30), Y(31), N0_31_61);
	-- signal N0_31_62 : std_logic;
	PP1675 : and2 port map (X(31), Y(31), N0_31_62);
	-- signal N0_31_63 : std_logic;
	PP1676 : and2 port map (X(32), Y(31), N0_31_63);
	-- signal N0_31_64 : std_logic;
	PP1677 : and2 port map (X(33), Y(31), N0_31_64);
	-- signal N0_31_65 : std_logic;
	PP1678 : and2 port map (X(34), Y(31), N0_31_65);
	-- signal N0_31_66 : std_logic;
	PP1679 : and2 port map (X(35), Y(31), N0_31_66);
	-- signal N0_31_67 : std_logic;
	PP1680 : and2 port map (X(36), Y(31), N0_31_67);
	-- signal N0_31_68 : std_logic;
	PP1681 : and2 port map (X(37), Y(31), N0_31_68);
	-- signal N0_31_69 : std_logic;
	PP1682 : and2 port map (X(38), Y(31), N0_31_69);
	-- signal N0_31_70 : std_logic;
	PP1683 : and2 port map (X(39), Y(31), N0_31_70);
	-- signal N0_31_71 : std_logic;
	PP1684 : and2 port map (X(40), Y(31), N0_31_71);
	-- signal N0_31_72 : std_logic;
	PP1685 : and2 port map (X(41), Y(31), N0_31_72);
	-- signal N0_31_73 : std_logic;
	PP1686 : and2 port map (X(42), Y(31), N0_31_73);
	-- signal N0_31_74 : std_logic;
	PP1687 : and2 port map (X(43), Y(31), N0_31_74);
	-- signal N0_31_75 : std_logic;
	PP1688 : and2 port map (X(44), Y(31), N0_31_75);
	-- signal N0_31_76 : std_logic;
	PP1689 : and2 port map (X(45), Y(31), N0_31_76);
	-- signal N0_31_77 : std_logic;
	PP1690 : and2 port map (X(46), Y(31), N0_31_77);
	-- signal N0_31_78 : std_logic;
	PP1691 : and2 port map (X(47), Y(31), N0_31_78);
	-- signal N0_31_79 : std_logic;
	PP1692 : and2 port map (X(48), Y(31), N0_31_79);
	-- signal N0_31_80 : std_logic;
	PP1693 : and2 port map (X(49), Y(31), N0_31_80);
	-- signal N0_31_81 : std_logic;
	PP1694 : and2 port map (X(50), Y(31), N0_31_81);
	-- signal N0_31_82 : std_logic;
	PP1695 : and2 port map (X(51), Y(31), N0_31_82);
	-- signal N0_31_83 : std_logic;
	PP1696 : and2 port map ('1', Y(31), N0_31_83);
	-- signal N0_32_32 : std_logic;
	PP1697 : and2 port map (X(0), Y(32), N0_32_32);
	-- signal N0_32_33 : std_logic;
	PP1698 : and2 port map (X(1), Y(32), N0_32_33);
	-- signal N0_32_34 : std_logic;
	PP1699 : and2 port map (X(2), Y(32), N0_32_34);
	-- signal N0_32_35 : std_logic;
	PP1700 : and2 port map (X(3), Y(32), N0_32_35);
	-- signal N0_32_36 : std_logic;
	PP1701 : and2 port map (X(4), Y(32), N0_32_36);
	-- signal N0_32_37 : std_logic;
	PP1702 : and2 port map (X(5), Y(32), N0_32_37);
	-- signal N0_32_38 : std_logic;
	PP1703 : and2 port map (X(6), Y(32), N0_32_38);
	-- signal N0_32_39 : std_logic;
	PP1704 : and2 port map (X(7), Y(32), N0_32_39);
	-- signal N0_32_40 : std_logic;
	PP1705 : and2 port map (X(8), Y(32), N0_32_40);
	-- signal N0_32_41 : std_logic;
	PP1706 : and2 port map (X(9), Y(32), N0_32_41);
	-- signal N0_32_42 : std_logic;
	PP1707 : and2 port map (X(10), Y(32), N0_32_42);
	-- signal N0_32_43 : std_logic;
	PP1708 : and2 port map (X(11), Y(32), N0_32_43);
	-- signal N0_32_44 : std_logic;
	PP1709 : and2 port map (X(12), Y(32), N0_32_44);
	-- signal N0_32_45 : std_logic;
	PP1710 : and2 port map (X(13), Y(32), N0_32_45);
	-- signal N0_32_46 : std_logic;
	PP1711 : and2 port map (X(14), Y(32), N0_32_46);
	-- signal N0_32_47 : std_logic;
	PP1712 : and2 port map (X(15), Y(32), N0_32_47);
	-- signal N0_32_48 : std_logic;
	PP1713 : and2 port map (X(16), Y(32), N0_32_48);
	-- signal N0_32_49 : std_logic;
	PP1714 : and2 port map (X(17), Y(32), N0_32_49);
	-- signal N0_32_50 : std_logic;
	PP1715 : and2 port map (X(18), Y(32), N0_32_50);
	-- signal N0_32_51 : std_logic;
	PP1716 : and2 port map (X(19), Y(32), N0_32_51);
	-- signal N0_32_52 : std_logic;
	PP1717 : and2 port map (X(20), Y(32), N0_32_52);
	-- signal N0_32_53 : std_logic;
	PP1718 : and2 port map (X(21), Y(32), N0_32_53);
	-- signal N0_32_54 : std_logic;
	PP1719 : and2 port map (X(22), Y(32), N0_32_54);
	-- signal N0_32_55 : std_logic;
	PP1720 : and2 port map (X(23), Y(32), N0_32_55);
	-- signal N0_32_56 : std_logic;
	PP1721 : and2 port map (X(24), Y(32), N0_32_56);
	-- signal N0_32_57 : std_logic;
	PP1722 : and2 port map (X(25), Y(32), N0_32_57);
	-- signal N0_32_58 : std_logic;
	PP1723 : and2 port map (X(26), Y(32), N0_32_58);
	-- signal N0_32_59 : std_logic;
	PP1724 : and2 port map (X(27), Y(32), N0_32_59);
	-- signal N0_32_60 : std_logic;
	PP1725 : and2 port map (X(28), Y(32), N0_32_60);
	-- signal N0_32_61 : std_logic;
	PP1726 : and2 port map (X(29), Y(32), N0_32_61);
	-- signal N0_32_62 : std_logic;
	PP1727 : and2 port map (X(30), Y(32), N0_32_62);
	-- signal N0_32_63 : std_logic;
	PP1728 : and2 port map (X(31), Y(32), N0_32_63);
	-- signal N0_32_64 : std_logic;
	PP1729 : and2 port map (X(32), Y(32), N0_32_64);
	-- signal N0_32_65 : std_logic;
	PP1730 : and2 port map (X(33), Y(32), N0_32_65);
	-- signal N0_32_66 : std_logic;
	PP1731 : and2 port map (X(34), Y(32), N0_32_66);
	-- signal N0_32_67 : std_logic;
	PP1732 : and2 port map (X(35), Y(32), N0_32_67);
	-- signal N0_32_68 : std_logic;
	PP1733 : and2 port map (X(36), Y(32), N0_32_68);
	-- signal N0_32_69 : std_logic;
	PP1734 : and2 port map (X(37), Y(32), N0_32_69);
	-- signal N0_32_70 : std_logic;
	PP1735 : and2 port map (X(38), Y(32), N0_32_70);
	-- signal N0_32_71 : std_logic;
	PP1736 : and2 port map (X(39), Y(32), N0_32_71);
	-- signal N0_32_72 : std_logic;
	PP1737 : and2 port map (X(40), Y(32), N0_32_72);
	-- signal N0_32_73 : std_logic;
	PP1738 : and2 port map (X(41), Y(32), N0_32_73);
	-- signal N0_32_74 : std_logic;
	PP1739 : and2 port map (X(42), Y(32), N0_32_74);
	-- signal N0_32_75 : std_logic;
	PP1740 : and2 port map (X(43), Y(32), N0_32_75);
	-- signal N0_32_76 : std_logic;
	PP1741 : and2 port map (X(44), Y(32), N0_32_76);
	-- signal N0_32_77 : std_logic;
	PP1742 : and2 port map (X(45), Y(32), N0_32_77);
	-- signal N0_32_78 : std_logic;
	PP1743 : and2 port map (X(46), Y(32), N0_32_78);
	-- signal N0_32_79 : std_logic;
	PP1744 : and2 port map (X(47), Y(32), N0_32_79);
	-- signal N0_32_80 : std_logic;
	PP1745 : and2 port map (X(48), Y(32), N0_32_80);
	-- signal N0_32_81 : std_logic;
	PP1746 : and2 port map (X(49), Y(32), N0_32_81);
	-- signal N0_32_82 : std_logic;
	PP1747 : and2 port map (X(50), Y(32), N0_32_82);
	-- signal N0_32_83 : std_logic;
	PP1748 : and2 port map (X(51), Y(32), N0_32_83);
	-- signal N0_32_84 : std_logic;
	PP1749 : and2 port map ('1', Y(32), N0_32_84);
	-- signal N0_33_33 : std_logic;
	PP1750 : and2 port map (X(0), Y(33), N0_33_33);
	-- signal N0_33_34 : std_logic;
	PP1751 : and2 port map (X(1), Y(33), N0_33_34);
	-- signal N0_33_35 : std_logic;
	PP1752 : and2 port map (X(2), Y(33), N0_33_35);
	-- signal N0_33_36 : std_logic;
	PP1753 : and2 port map (X(3), Y(33), N0_33_36);
	-- signal N0_33_37 : std_logic;
	PP1754 : and2 port map (X(4), Y(33), N0_33_37);
	-- signal N0_33_38 : std_logic;
	PP1755 : and2 port map (X(5), Y(33), N0_33_38);
	-- signal N0_33_39 : std_logic;
	PP1756 : and2 port map (X(6), Y(33), N0_33_39);
	-- signal N0_33_40 : std_logic;
	PP1757 : and2 port map (X(7), Y(33), N0_33_40);
	-- signal N0_33_41 : std_logic;
	PP1758 : and2 port map (X(8), Y(33), N0_33_41);
	-- signal N0_33_42 : std_logic;
	PP1759 : and2 port map (X(9), Y(33), N0_33_42);
	-- signal N0_33_43 : std_logic;
	PP1760 : and2 port map (X(10), Y(33), N0_33_43);
	-- signal N0_33_44 : std_logic;
	PP1761 : and2 port map (X(11), Y(33), N0_33_44);
	-- signal N0_33_45 : std_logic;
	PP1762 : and2 port map (X(12), Y(33), N0_33_45);
	-- signal N0_33_46 : std_logic;
	PP1763 : and2 port map (X(13), Y(33), N0_33_46);
	-- signal N0_33_47 : std_logic;
	PP1764 : and2 port map (X(14), Y(33), N0_33_47);
	-- signal N0_33_48 : std_logic;
	PP1765 : and2 port map (X(15), Y(33), N0_33_48);
	-- signal N0_33_49 : std_logic;
	PP1766 : and2 port map (X(16), Y(33), N0_33_49);
	-- signal N0_33_50 : std_logic;
	PP1767 : and2 port map (X(17), Y(33), N0_33_50);
	-- signal N0_33_51 : std_logic;
	PP1768 : and2 port map (X(18), Y(33), N0_33_51);
	-- signal N0_33_52 : std_logic;
	PP1769 : and2 port map (X(19), Y(33), N0_33_52);
	-- signal N0_33_53 : std_logic;
	PP1770 : and2 port map (X(20), Y(33), N0_33_53);
	-- signal N0_33_54 : std_logic;
	PP1771 : and2 port map (X(21), Y(33), N0_33_54);
	-- signal N0_33_55 : std_logic;
	PP1772 : and2 port map (X(22), Y(33), N0_33_55);
	-- signal N0_33_56 : std_logic;
	PP1773 : and2 port map (X(23), Y(33), N0_33_56);
	-- signal N0_33_57 : std_logic;
	PP1774 : and2 port map (X(24), Y(33), N0_33_57);
	-- signal N0_33_58 : std_logic;
	PP1775 : and2 port map (X(25), Y(33), N0_33_58);
	-- signal N0_33_59 : std_logic;
	PP1776 : and2 port map (X(26), Y(33), N0_33_59);
	-- signal N0_33_60 : std_logic;
	PP1777 : and2 port map (X(27), Y(33), N0_33_60);
	-- signal N0_33_61 : std_logic;
	PP1778 : and2 port map (X(28), Y(33), N0_33_61);
	-- signal N0_33_62 : std_logic;
	PP1779 : and2 port map (X(29), Y(33), N0_33_62);
	-- signal N0_33_63 : std_logic;
	PP1780 : and2 port map (X(30), Y(33), N0_33_63);
	-- signal N0_33_64 : std_logic;
	PP1781 : and2 port map (X(31), Y(33), N0_33_64);
	-- signal N0_33_65 : std_logic;
	PP1782 : and2 port map (X(32), Y(33), N0_33_65);
	-- signal N0_33_66 : std_logic;
	PP1783 : and2 port map (X(33), Y(33), N0_33_66);
	-- signal N0_33_67 : std_logic;
	PP1784 : and2 port map (X(34), Y(33), N0_33_67);
	-- signal N0_33_68 : std_logic;
	PP1785 : and2 port map (X(35), Y(33), N0_33_68);
	-- signal N0_33_69 : std_logic;
	PP1786 : and2 port map (X(36), Y(33), N0_33_69);
	-- signal N0_33_70 : std_logic;
	PP1787 : and2 port map (X(37), Y(33), N0_33_70);
	-- signal N0_33_71 : std_logic;
	PP1788 : and2 port map (X(38), Y(33), N0_33_71);
	-- signal N0_33_72 : std_logic;
	PP1789 : and2 port map (X(39), Y(33), N0_33_72);
	-- signal N0_33_73 : std_logic;
	PP1790 : and2 port map (X(40), Y(33), N0_33_73);
	-- signal N0_33_74 : std_logic;
	PP1791 : and2 port map (X(41), Y(33), N0_33_74);
	-- signal N0_33_75 : std_logic;
	PP1792 : and2 port map (X(42), Y(33), N0_33_75);
	-- signal N0_33_76 : std_logic;
	PP1793 : and2 port map (X(43), Y(33), N0_33_76);
	-- signal N0_33_77 : std_logic;
	PP1794 : and2 port map (X(44), Y(33), N0_33_77);
	-- signal N0_33_78 : std_logic;
	PP1795 : and2 port map (X(45), Y(33), N0_33_78);
	-- signal N0_33_79 : std_logic;
	PP1796 : and2 port map (X(46), Y(33), N0_33_79);
	-- signal N0_33_80 : std_logic;
	PP1797 : and2 port map (X(47), Y(33), N0_33_80);
	-- signal N0_33_81 : std_logic;
	PP1798 : and2 port map (X(48), Y(33), N0_33_81);
	-- signal N0_33_82 : std_logic;
	PP1799 : and2 port map (X(49), Y(33), N0_33_82);
	-- signal N0_33_83 : std_logic;
	PP1800 : and2 port map (X(50), Y(33), N0_33_83);
	-- signal N0_33_84 : std_logic;
	PP1801 : and2 port map (X(51), Y(33), N0_33_84);
	-- signal N0_33_85 : std_logic;
	PP1802 : and2 port map ('1', Y(33), N0_33_85);
	-- signal N0_34_34 : std_logic;
	PP1803 : and2 port map (X(0), Y(34), N0_34_34);
	-- signal N0_34_35 : std_logic;
	PP1804 : and2 port map (X(1), Y(34), N0_34_35);
	-- signal N0_34_36 : std_logic;
	PP1805 : and2 port map (X(2), Y(34), N0_34_36);
	-- signal N0_34_37 : std_logic;
	PP1806 : and2 port map (X(3), Y(34), N0_34_37);
	-- signal N0_34_38 : std_logic;
	PP1807 : and2 port map (X(4), Y(34), N0_34_38);
	-- signal N0_34_39 : std_logic;
	PP1808 : and2 port map (X(5), Y(34), N0_34_39);
	-- signal N0_34_40 : std_logic;
	PP1809 : and2 port map (X(6), Y(34), N0_34_40);
	-- signal N0_34_41 : std_logic;
	PP1810 : and2 port map (X(7), Y(34), N0_34_41);
	-- signal N0_34_42 : std_logic;
	PP1811 : and2 port map (X(8), Y(34), N0_34_42);
	-- signal N0_34_43 : std_logic;
	PP1812 : and2 port map (X(9), Y(34), N0_34_43);
	-- signal N0_34_44 : std_logic;
	PP1813 : and2 port map (X(10), Y(34), N0_34_44);
	-- signal N0_34_45 : std_logic;
	PP1814 : and2 port map (X(11), Y(34), N0_34_45);
	-- signal N0_34_46 : std_logic;
	PP1815 : and2 port map (X(12), Y(34), N0_34_46);
	-- signal N0_34_47 : std_logic;
	PP1816 : and2 port map (X(13), Y(34), N0_34_47);
	-- signal N0_34_48 : std_logic;
	PP1817 : and2 port map (X(14), Y(34), N0_34_48);
	-- signal N0_34_49 : std_logic;
	PP1818 : and2 port map (X(15), Y(34), N0_34_49);
	-- signal N0_34_50 : std_logic;
	PP1819 : and2 port map (X(16), Y(34), N0_34_50);
	-- signal N0_34_51 : std_logic;
	PP1820 : and2 port map (X(17), Y(34), N0_34_51);
	-- signal N0_34_52 : std_logic;
	PP1821 : and2 port map (X(18), Y(34), N0_34_52);
	-- signal N0_34_53 : std_logic;
	PP1822 : and2 port map (X(19), Y(34), N0_34_53);
	-- signal N0_34_54 : std_logic;
	PP1823 : and2 port map (X(20), Y(34), N0_34_54);
	-- signal N0_34_55 : std_logic;
	PP1824 : and2 port map (X(21), Y(34), N0_34_55);
	-- signal N0_34_56 : std_logic;
	PP1825 : and2 port map (X(22), Y(34), N0_34_56);
	-- signal N0_34_57 : std_logic;
	PP1826 : and2 port map (X(23), Y(34), N0_34_57);
	-- signal N0_34_58 : std_logic;
	PP1827 : and2 port map (X(24), Y(34), N0_34_58);
	-- signal N0_34_59 : std_logic;
	PP1828 : and2 port map (X(25), Y(34), N0_34_59);
	-- signal N0_34_60 : std_logic;
	PP1829 : and2 port map (X(26), Y(34), N0_34_60);
	-- signal N0_34_61 : std_logic;
	PP1830 : and2 port map (X(27), Y(34), N0_34_61);
	-- signal N0_34_62 : std_logic;
	PP1831 : and2 port map (X(28), Y(34), N0_34_62);
	-- signal N0_34_63 : std_logic;
	PP1832 : and2 port map (X(29), Y(34), N0_34_63);
	-- signal N0_34_64 : std_logic;
	PP1833 : and2 port map (X(30), Y(34), N0_34_64);
	-- signal N0_34_65 : std_logic;
	PP1834 : and2 port map (X(31), Y(34), N0_34_65);
	-- signal N0_34_66 : std_logic;
	PP1835 : and2 port map (X(32), Y(34), N0_34_66);
	-- signal N0_34_67 : std_logic;
	PP1836 : and2 port map (X(33), Y(34), N0_34_67);
	-- signal N0_34_68 : std_logic;
	PP1837 : and2 port map (X(34), Y(34), N0_34_68);
	-- signal N0_34_69 : std_logic;
	PP1838 : and2 port map (X(35), Y(34), N0_34_69);
	-- signal N0_34_70 : std_logic;
	PP1839 : and2 port map (X(36), Y(34), N0_34_70);
	-- signal N0_34_71 : std_logic;
	PP1840 : and2 port map (X(37), Y(34), N0_34_71);
	-- signal N0_34_72 : std_logic;
	PP1841 : and2 port map (X(38), Y(34), N0_34_72);
	-- signal N0_34_73 : std_logic;
	PP1842 : and2 port map (X(39), Y(34), N0_34_73);
	-- signal N0_34_74 : std_logic;
	PP1843 : and2 port map (X(40), Y(34), N0_34_74);
	-- signal N0_34_75 : std_logic;
	PP1844 : and2 port map (X(41), Y(34), N0_34_75);
	-- signal N0_34_76 : std_logic;
	PP1845 : and2 port map (X(42), Y(34), N0_34_76);
	-- signal N0_34_77 : std_logic;
	PP1846 : and2 port map (X(43), Y(34), N0_34_77);
	-- signal N0_34_78 : std_logic;
	PP1847 : and2 port map (X(44), Y(34), N0_34_78);
	-- signal N0_34_79 : std_logic;
	PP1848 : and2 port map (X(45), Y(34), N0_34_79);
	-- signal N0_34_80 : std_logic;
	PP1849 : and2 port map (X(46), Y(34), N0_34_80);
	-- signal N0_34_81 : std_logic;
	PP1850 : and2 port map (X(47), Y(34), N0_34_81);
	-- signal N0_34_82 : std_logic;
	PP1851 : and2 port map (X(48), Y(34), N0_34_82);
	-- signal N0_34_83 : std_logic;
	PP1852 : and2 port map (X(49), Y(34), N0_34_83);
	-- signal N0_34_84 : std_logic;
	PP1853 : and2 port map (X(50), Y(34), N0_34_84);
	-- signal N0_34_85 : std_logic;
	PP1854 : and2 port map (X(51), Y(34), N0_34_85);
	-- signal N0_34_86 : std_logic;
	PP1855 : and2 port map ('1', Y(34), N0_34_86);
	-- signal N0_35_35 : std_logic;
	PP1856 : and2 port map (X(0), Y(35), N0_35_35);
	-- signal N0_35_36 : std_logic;
	PP1857 : and2 port map (X(1), Y(35), N0_35_36);
	-- signal N0_35_37 : std_logic;
	PP1858 : and2 port map (X(2), Y(35), N0_35_37);
	-- signal N0_35_38 : std_logic;
	PP1859 : and2 port map (X(3), Y(35), N0_35_38);
	-- signal N0_35_39 : std_logic;
	PP1860 : and2 port map (X(4), Y(35), N0_35_39);
	-- signal N0_35_40 : std_logic;
	PP1861 : and2 port map (X(5), Y(35), N0_35_40);
	-- signal N0_35_41 : std_logic;
	PP1862 : and2 port map (X(6), Y(35), N0_35_41);
	-- signal N0_35_42 : std_logic;
	PP1863 : and2 port map (X(7), Y(35), N0_35_42);
	-- signal N0_35_43 : std_logic;
	PP1864 : and2 port map (X(8), Y(35), N0_35_43);
	-- signal N0_35_44 : std_logic;
	PP1865 : and2 port map (X(9), Y(35), N0_35_44);
	-- signal N0_35_45 : std_logic;
	PP1866 : and2 port map (X(10), Y(35), N0_35_45);
	-- signal N0_35_46 : std_logic;
	PP1867 : and2 port map (X(11), Y(35), N0_35_46);
	-- signal N0_35_47 : std_logic;
	PP1868 : and2 port map (X(12), Y(35), N0_35_47);
	-- signal N0_35_48 : std_logic;
	PP1869 : and2 port map (X(13), Y(35), N0_35_48);
	-- signal N0_35_49 : std_logic;
	PP1870 : and2 port map (X(14), Y(35), N0_35_49);
	-- signal N0_35_50 : std_logic;
	PP1871 : and2 port map (X(15), Y(35), N0_35_50);
	-- signal N0_35_51 : std_logic;
	PP1872 : and2 port map (X(16), Y(35), N0_35_51);
	-- signal N0_35_52 : std_logic;
	PP1873 : and2 port map (X(17), Y(35), N0_35_52);
	-- signal N0_35_53 : std_logic;
	PP1874 : and2 port map (X(18), Y(35), N0_35_53);
	-- signal N0_35_54 : std_logic;
	PP1875 : and2 port map (X(19), Y(35), N0_35_54);
	-- signal N0_35_55 : std_logic;
	PP1876 : and2 port map (X(20), Y(35), N0_35_55);
	-- signal N0_35_56 : std_logic;
	PP1877 : and2 port map (X(21), Y(35), N0_35_56);
	-- signal N0_35_57 : std_logic;
	PP1878 : and2 port map (X(22), Y(35), N0_35_57);
	-- signal N0_35_58 : std_logic;
	PP1879 : and2 port map (X(23), Y(35), N0_35_58);
	-- signal N0_35_59 : std_logic;
	PP1880 : and2 port map (X(24), Y(35), N0_35_59);
	-- signal N0_35_60 : std_logic;
	PP1881 : and2 port map (X(25), Y(35), N0_35_60);
	-- signal N0_35_61 : std_logic;
	PP1882 : and2 port map (X(26), Y(35), N0_35_61);
	-- signal N0_35_62 : std_logic;
	PP1883 : and2 port map (X(27), Y(35), N0_35_62);
	-- signal N0_35_63 : std_logic;
	PP1884 : and2 port map (X(28), Y(35), N0_35_63);
	-- signal N0_35_64 : std_logic;
	PP1885 : and2 port map (X(29), Y(35), N0_35_64);
	-- signal N0_35_65 : std_logic;
	PP1886 : and2 port map (X(30), Y(35), N0_35_65);
	-- signal N0_35_66 : std_logic;
	PP1887 : and2 port map (X(31), Y(35), N0_35_66);
	-- signal N0_35_67 : std_logic;
	PP1888 : and2 port map (X(32), Y(35), N0_35_67);
	-- signal N0_35_68 : std_logic;
	PP1889 : and2 port map (X(33), Y(35), N0_35_68);
	-- signal N0_35_69 : std_logic;
	PP1890 : and2 port map (X(34), Y(35), N0_35_69);
	-- signal N0_35_70 : std_logic;
	PP1891 : and2 port map (X(35), Y(35), N0_35_70);
	-- signal N0_35_71 : std_logic;
	PP1892 : and2 port map (X(36), Y(35), N0_35_71);
	-- signal N0_35_72 : std_logic;
	PP1893 : and2 port map (X(37), Y(35), N0_35_72);
	-- signal N0_35_73 : std_logic;
	PP1894 : and2 port map (X(38), Y(35), N0_35_73);
	-- signal N0_35_74 : std_logic;
	PP1895 : and2 port map (X(39), Y(35), N0_35_74);
	-- signal N0_35_75 : std_logic;
	PP1896 : and2 port map (X(40), Y(35), N0_35_75);
	-- signal N0_35_76 : std_logic;
	PP1897 : and2 port map (X(41), Y(35), N0_35_76);
	-- signal N0_35_77 : std_logic;
	PP1898 : and2 port map (X(42), Y(35), N0_35_77);
	-- signal N0_35_78 : std_logic;
	PP1899 : and2 port map (X(43), Y(35), N0_35_78);
	-- signal N0_35_79 : std_logic;
	PP1900 : and2 port map (X(44), Y(35), N0_35_79);
	-- signal N0_35_80 : std_logic;
	PP1901 : and2 port map (X(45), Y(35), N0_35_80);
	-- signal N0_35_81 : std_logic;
	PP1902 : and2 port map (X(46), Y(35), N0_35_81);
	-- signal N0_35_82 : std_logic;
	PP1903 : and2 port map (X(47), Y(35), N0_35_82);
	-- signal N0_35_83 : std_logic;
	PP1904 : and2 port map (X(48), Y(35), N0_35_83);
	-- signal N0_35_84 : std_logic;
	PP1905 : and2 port map (X(49), Y(35), N0_35_84);
	-- signal N0_35_85 : std_logic;
	PP1906 : and2 port map (X(50), Y(35), N0_35_85);
	-- signal N0_35_86 : std_logic;
	PP1907 : and2 port map (X(51), Y(35), N0_35_86);
	-- signal N0_35_87 : std_logic;
	PP1908 : and2 port map ('1', Y(35), N0_35_87);
	-- signal N0_36_36 : std_logic;
	PP1909 : and2 port map (X(0), Y(36), N0_36_36);
	-- signal N0_36_37 : std_logic;
	PP1910 : and2 port map (X(1), Y(36), N0_36_37);
	-- signal N0_36_38 : std_logic;
	PP1911 : and2 port map (X(2), Y(36), N0_36_38);
	-- signal N0_36_39 : std_logic;
	PP1912 : and2 port map (X(3), Y(36), N0_36_39);
	-- signal N0_36_40 : std_logic;
	PP1913 : and2 port map (X(4), Y(36), N0_36_40);
	-- signal N0_36_41 : std_logic;
	PP1914 : and2 port map (X(5), Y(36), N0_36_41);
	-- signal N0_36_42 : std_logic;
	PP1915 : and2 port map (X(6), Y(36), N0_36_42);
	-- signal N0_36_43 : std_logic;
	PP1916 : and2 port map (X(7), Y(36), N0_36_43);
	-- signal N0_36_44 : std_logic;
	PP1917 : and2 port map (X(8), Y(36), N0_36_44);
	-- signal N0_36_45 : std_logic;
	PP1918 : and2 port map (X(9), Y(36), N0_36_45);
	-- signal N0_36_46 : std_logic;
	PP1919 : and2 port map (X(10), Y(36), N0_36_46);
	-- signal N0_36_47 : std_logic;
	PP1920 : and2 port map (X(11), Y(36), N0_36_47);
	-- signal N0_36_48 : std_logic;
	PP1921 : and2 port map (X(12), Y(36), N0_36_48);
	-- signal N0_36_49 : std_logic;
	PP1922 : and2 port map (X(13), Y(36), N0_36_49);
	-- signal N0_36_50 : std_logic;
	PP1923 : and2 port map (X(14), Y(36), N0_36_50);
	-- signal N0_36_51 : std_logic;
	PP1924 : and2 port map (X(15), Y(36), N0_36_51);
	-- signal N0_36_52 : std_logic;
	PP1925 : and2 port map (X(16), Y(36), N0_36_52);
	-- signal N0_36_53 : std_logic;
	PP1926 : and2 port map (X(17), Y(36), N0_36_53);
	-- signal N0_36_54 : std_logic;
	PP1927 : and2 port map (X(18), Y(36), N0_36_54);
	-- signal N0_36_55 : std_logic;
	PP1928 : and2 port map (X(19), Y(36), N0_36_55);
	-- signal N0_36_56 : std_logic;
	PP1929 : and2 port map (X(20), Y(36), N0_36_56);
	-- signal N0_36_57 : std_logic;
	PP1930 : and2 port map (X(21), Y(36), N0_36_57);
	-- signal N0_36_58 : std_logic;
	PP1931 : and2 port map (X(22), Y(36), N0_36_58);
	-- signal N0_36_59 : std_logic;
	PP1932 : and2 port map (X(23), Y(36), N0_36_59);
	-- signal N0_36_60 : std_logic;
	PP1933 : and2 port map (X(24), Y(36), N0_36_60);
	-- signal N0_36_61 : std_logic;
	PP1934 : and2 port map (X(25), Y(36), N0_36_61);
	-- signal N0_36_62 : std_logic;
	PP1935 : and2 port map (X(26), Y(36), N0_36_62);
	-- signal N0_36_63 : std_logic;
	PP1936 : and2 port map (X(27), Y(36), N0_36_63);
	-- signal N0_36_64 : std_logic;
	PP1937 : and2 port map (X(28), Y(36), N0_36_64);
	-- signal N0_36_65 : std_logic;
	PP1938 : and2 port map (X(29), Y(36), N0_36_65);
	-- signal N0_36_66 : std_logic;
	PP1939 : and2 port map (X(30), Y(36), N0_36_66);
	-- signal N0_36_67 : std_logic;
	PP1940 : and2 port map (X(31), Y(36), N0_36_67);
	-- signal N0_36_68 : std_logic;
	PP1941 : and2 port map (X(32), Y(36), N0_36_68);
	-- signal N0_36_69 : std_logic;
	PP1942 : and2 port map (X(33), Y(36), N0_36_69);
	-- signal N0_36_70 : std_logic;
	PP1943 : and2 port map (X(34), Y(36), N0_36_70);
	-- signal N0_36_71 : std_logic;
	PP1944 : and2 port map (X(35), Y(36), N0_36_71);
	-- signal N0_36_72 : std_logic;
	PP1945 : and2 port map (X(36), Y(36), N0_36_72);
	-- signal N0_36_73 : std_logic;
	PP1946 : and2 port map (X(37), Y(36), N0_36_73);
	-- signal N0_36_74 : std_logic;
	PP1947 : and2 port map (X(38), Y(36), N0_36_74);
	-- signal N0_36_75 : std_logic;
	PP1948 : and2 port map (X(39), Y(36), N0_36_75);
	-- signal N0_36_76 : std_logic;
	PP1949 : and2 port map (X(40), Y(36), N0_36_76);
	-- signal N0_36_77 : std_logic;
	PP1950 : and2 port map (X(41), Y(36), N0_36_77);
	-- signal N0_36_78 : std_logic;
	PP1951 : and2 port map (X(42), Y(36), N0_36_78);
	-- signal N0_36_79 : std_logic;
	PP1952 : and2 port map (X(43), Y(36), N0_36_79);
	-- signal N0_36_80 : std_logic;
	PP1953 : and2 port map (X(44), Y(36), N0_36_80);
	-- signal N0_36_81 : std_logic;
	PP1954 : and2 port map (X(45), Y(36), N0_36_81);
	-- signal N0_36_82 : std_logic;
	PP1955 : and2 port map (X(46), Y(36), N0_36_82);
	-- signal N0_36_83 : std_logic;
	PP1956 : and2 port map (X(47), Y(36), N0_36_83);
	-- signal N0_36_84 : std_logic;
	PP1957 : and2 port map (X(48), Y(36), N0_36_84);
	-- signal N0_36_85 : std_logic;
	PP1958 : and2 port map (X(49), Y(36), N0_36_85);
	-- signal N0_36_86 : std_logic;
	PP1959 : and2 port map (X(50), Y(36), N0_36_86);
	-- signal N0_36_87 : std_logic;
	PP1960 : and2 port map (X(51), Y(36), N0_36_87);
	-- signal N0_36_88 : std_logic;
	PP1961 : and2 port map ('1', Y(36), N0_36_88);
	-- signal N0_37_37 : std_logic;
	PP1962 : and2 port map (X(0), Y(37), N0_37_37);
	-- signal N0_37_38 : std_logic;
	PP1963 : and2 port map (X(1), Y(37), N0_37_38);
	-- signal N0_37_39 : std_logic;
	PP1964 : and2 port map (X(2), Y(37), N0_37_39);
	-- signal N0_37_40 : std_logic;
	PP1965 : and2 port map (X(3), Y(37), N0_37_40);
	-- signal N0_37_41 : std_logic;
	PP1966 : and2 port map (X(4), Y(37), N0_37_41);
	-- signal N0_37_42 : std_logic;
	PP1967 : and2 port map (X(5), Y(37), N0_37_42);
	-- signal N0_37_43 : std_logic;
	PP1968 : and2 port map (X(6), Y(37), N0_37_43);
	-- signal N0_37_44 : std_logic;
	PP1969 : and2 port map (X(7), Y(37), N0_37_44);
	-- signal N0_37_45 : std_logic;
	PP1970 : and2 port map (X(8), Y(37), N0_37_45);
	-- signal N0_37_46 : std_logic;
	PP1971 : and2 port map (X(9), Y(37), N0_37_46);
	-- signal N0_37_47 : std_logic;
	PP1972 : and2 port map (X(10), Y(37), N0_37_47);
	-- signal N0_37_48 : std_logic;
	PP1973 : and2 port map (X(11), Y(37), N0_37_48);
	-- signal N0_37_49 : std_logic;
	PP1974 : and2 port map (X(12), Y(37), N0_37_49);
	-- signal N0_37_50 : std_logic;
	PP1975 : and2 port map (X(13), Y(37), N0_37_50);
	-- signal N0_37_51 : std_logic;
	PP1976 : and2 port map (X(14), Y(37), N0_37_51);
	-- signal N0_37_52 : std_logic;
	PP1977 : and2 port map (X(15), Y(37), N0_37_52);
	-- signal N0_37_53 : std_logic;
	PP1978 : and2 port map (X(16), Y(37), N0_37_53);
	-- signal N0_37_54 : std_logic;
	PP1979 : and2 port map (X(17), Y(37), N0_37_54);
	-- signal N0_37_55 : std_logic;
	PP1980 : and2 port map (X(18), Y(37), N0_37_55);
	-- signal N0_37_56 : std_logic;
	PP1981 : and2 port map (X(19), Y(37), N0_37_56);
	-- signal N0_37_57 : std_logic;
	PP1982 : and2 port map (X(20), Y(37), N0_37_57);
	-- signal N0_37_58 : std_logic;
	PP1983 : and2 port map (X(21), Y(37), N0_37_58);
	-- signal N0_37_59 : std_logic;
	PP1984 : and2 port map (X(22), Y(37), N0_37_59);
	-- signal N0_37_60 : std_logic;
	PP1985 : and2 port map (X(23), Y(37), N0_37_60);
	-- signal N0_37_61 : std_logic;
	PP1986 : and2 port map (X(24), Y(37), N0_37_61);
	-- signal N0_37_62 : std_logic;
	PP1987 : and2 port map (X(25), Y(37), N0_37_62);
	-- signal N0_37_63 : std_logic;
	PP1988 : and2 port map (X(26), Y(37), N0_37_63);
	-- signal N0_37_64 : std_logic;
	PP1989 : and2 port map (X(27), Y(37), N0_37_64);
	-- signal N0_37_65 : std_logic;
	PP1990 : and2 port map (X(28), Y(37), N0_37_65);
	-- signal N0_37_66 : std_logic;
	PP1991 : and2 port map (X(29), Y(37), N0_37_66);
	-- signal N0_37_67 : std_logic;
	PP1992 : and2 port map (X(30), Y(37), N0_37_67);
	-- signal N0_37_68 : std_logic;
	PP1993 : and2 port map (X(31), Y(37), N0_37_68);
	-- signal N0_37_69 : std_logic;
	PP1994 : and2 port map (X(32), Y(37), N0_37_69);
	-- signal N0_37_70 : std_logic;
	PP1995 : and2 port map (X(33), Y(37), N0_37_70);
	-- signal N0_37_71 : std_logic;
	PP1996 : and2 port map (X(34), Y(37), N0_37_71);
	-- signal N0_37_72 : std_logic;
	PP1997 : and2 port map (X(35), Y(37), N0_37_72);
	-- signal N0_37_73 : std_logic;
	PP1998 : and2 port map (X(36), Y(37), N0_37_73);
	-- signal N0_37_74 : std_logic;
	PP1999 : and2 port map (X(37), Y(37), N0_37_74);
	-- signal N0_37_75 : std_logic;
	PP2000 : and2 port map (X(38), Y(37), N0_37_75);
	-- signal N0_37_76 : std_logic;
	PP2001 : and2 port map (X(39), Y(37), N0_37_76);
	-- signal N0_37_77 : std_logic;
	PP2002 : and2 port map (X(40), Y(37), N0_37_77);
	-- signal N0_37_78 : std_logic;
	PP2003 : and2 port map (X(41), Y(37), N0_37_78);
	-- signal N0_37_79 : std_logic;
	PP2004 : and2 port map (X(42), Y(37), N0_37_79);
	-- signal N0_37_80 : std_logic;
	PP2005 : and2 port map (X(43), Y(37), N0_37_80);
	-- signal N0_37_81 : std_logic;
	PP2006 : and2 port map (X(44), Y(37), N0_37_81);
	-- signal N0_37_82 : std_logic;
	PP2007 : and2 port map (X(45), Y(37), N0_37_82);
	-- signal N0_37_83 : std_logic;
	PP2008 : and2 port map (X(46), Y(37), N0_37_83);
	-- signal N0_37_84 : std_logic;
	PP2009 : and2 port map (X(47), Y(37), N0_37_84);
	-- signal N0_37_85 : std_logic;
	PP2010 : and2 port map (X(48), Y(37), N0_37_85);
	-- signal N0_37_86 : std_logic;
	PP2011 : and2 port map (X(49), Y(37), N0_37_86);
	-- signal N0_37_87 : std_logic;
	PP2012 : and2 port map (X(50), Y(37), N0_37_87);
	-- signal N0_37_88 : std_logic;
	PP2013 : and2 port map (X(51), Y(37), N0_37_88);
	-- signal N0_37_89 : std_logic;
	PP2014 : and2 port map ('1', Y(37), N0_37_89);
	-- signal N0_38_38 : std_logic;
	PP2015 : and2 port map (X(0), Y(38), N0_38_38);
	-- signal N0_38_39 : std_logic;
	PP2016 : and2 port map (X(1), Y(38), N0_38_39);
	-- signal N0_38_40 : std_logic;
	PP2017 : and2 port map (X(2), Y(38), N0_38_40);
	-- signal N0_38_41 : std_logic;
	PP2018 : and2 port map (X(3), Y(38), N0_38_41);
	-- signal N0_38_42 : std_logic;
	PP2019 : and2 port map (X(4), Y(38), N0_38_42);
	-- signal N0_38_43 : std_logic;
	PP2020 : and2 port map (X(5), Y(38), N0_38_43);
	-- signal N0_38_44 : std_logic;
	PP2021 : and2 port map (X(6), Y(38), N0_38_44);
	-- signal N0_38_45 : std_logic;
	PP2022 : and2 port map (X(7), Y(38), N0_38_45);
	-- signal N0_38_46 : std_logic;
	PP2023 : and2 port map (X(8), Y(38), N0_38_46);
	-- signal N0_38_47 : std_logic;
	PP2024 : and2 port map (X(9), Y(38), N0_38_47);
	-- signal N0_38_48 : std_logic;
	PP2025 : and2 port map (X(10), Y(38), N0_38_48);
	-- signal N0_38_49 : std_logic;
	PP2026 : and2 port map (X(11), Y(38), N0_38_49);
	-- signal N0_38_50 : std_logic;
	PP2027 : and2 port map (X(12), Y(38), N0_38_50);
	-- signal N0_38_51 : std_logic;
	PP2028 : and2 port map (X(13), Y(38), N0_38_51);
	-- signal N0_38_52 : std_logic;
	PP2029 : and2 port map (X(14), Y(38), N0_38_52);
	-- signal N0_38_53 : std_logic;
	PP2030 : and2 port map (X(15), Y(38), N0_38_53);
	-- signal N0_38_54 : std_logic;
	PP2031 : and2 port map (X(16), Y(38), N0_38_54);
	-- signal N0_38_55 : std_logic;
	PP2032 : and2 port map (X(17), Y(38), N0_38_55);
	-- signal N0_38_56 : std_logic;
	PP2033 : and2 port map (X(18), Y(38), N0_38_56);
	-- signal N0_38_57 : std_logic;
	PP2034 : and2 port map (X(19), Y(38), N0_38_57);
	-- signal N0_38_58 : std_logic;
	PP2035 : and2 port map (X(20), Y(38), N0_38_58);
	-- signal N0_38_59 : std_logic;
	PP2036 : and2 port map (X(21), Y(38), N0_38_59);
	-- signal N0_38_60 : std_logic;
	PP2037 : and2 port map (X(22), Y(38), N0_38_60);
	-- signal N0_38_61 : std_logic;
	PP2038 : and2 port map (X(23), Y(38), N0_38_61);
	-- signal N0_38_62 : std_logic;
	PP2039 : and2 port map (X(24), Y(38), N0_38_62);
	-- signal N0_38_63 : std_logic;
	PP2040 : and2 port map (X(25), Y(38), N0_38_63);
	-- signal N0_38_64 : std_logic;
	PP2041 : and2 port map (X(26), Y(38), N0_38_64);
	-- signal N0_38_65 : std_logic;
	PP2042 : and2 port map (X(27), Y(38), N0_38_65);
	-- signal N0_38_66 : std_logic;
	PP2043 : and2 port map (X(28), Y(38), N0_38_66);
	-- signal N0_38_67 : std_logic;
	PP2044 : and2 port map (X(29), Y(38), N0_38_67);
	-- signal N0_38_68 : std_logic;
	PP2045 : and2 port map (X(30), Y(38), N0_38_68);
	-- signal N0_38_69 : std_logic;
	PP2046 : and2 port map (X(31), Y(38), N0_38_69);
	-- signal N0_38_70 : std_logic;
	PP2047 : and2 port map (X(32), Y(38), N0_38_70);
	-- signal N0_38_71 : std_logic;
	PP2048 : and2 port map (X(33), Y(38), N0_38_71);
	-- signal N0_38_72 : std_logic;
	PP2049 : and2 port map (X(34), Y(38), N0_38_72);
	-- signal N0_38_73 : std_logic;
	PP2050 : and2 port map (X(35), Y(38), N0_38_73);
	-- signal N0_38_74 : std_logic;
	PP2051 : and2 port map (X(36), Y(38), N0_38_74);
	-- signal N0_38_75 : std_logic;
	PP2052 : and2 port map (X(37), Y(38), N0_38_75);
	-- signal N0_38_76 : std_logic;
	PP2053 : and2 port map (X(38), Y(38), N0_38_76);
	-- signal N0_38_77 : std_logic;
	PP2054 : and2 port map (X(39), Y(38), N0_38_77);
	-- signal N0_38_78 : std_logic;
	PP2055 : and2 port map (X(40), Y(38), N0_38_78);
	-- signal N0_38_79 : std_logic;
	PP2056 : and2 port map (X(41), Y(38), N0_38_79);
	-- signal N0_38_80 : std_logic;
	PP2057 : and2 port map (X(42), Y(38), N0_38_80);
	-- signal N0_38_81 : std_logic;
	PP2058 : and2 port map (X(43), Y(38), N0_38_81);
	-- signal N0_38_82 : std_logic;
	PP2059 : and2 port map (X(44), Y(38), N0_38_82);
	-- signal N0_38_83 : std_logic;
	PP2060 : and2 port map (X(45), Y(38), N0_38_83);
	-- signal N0_38_84 : std_logic;
	PP2061 : and2 port map (X(46), Y(38), N0_38_84);
	-- signal N0_38_85 : std_logic;
	PP2062 : and2 port map (X(47), Y(38), N0_38_85);
	-- signal N0_38_86 : std_logic;
	PP2063 : and2 port map (X(48), Y(38), N0_38_86);
	-- signal N0_38_87 : std_logic;
	PP2064 : and2 port map (X(49), Y(38), N0_38_87);
	-- signal N0_38_88 : std_logic;
	PP2065 : and2 port map (X(50), Y(38), N0_38_88);
	-- signal N0_38_89 : std_logic;
	PP2066 : and2 port map (X(51), Y(38), N0_38_89);
	-- signal N0_38_90 : std_logic;
	PP2067 : and2 port map ('1', Y(38), N0_38_90);
	-- signal N0_39_39 : std_logic;
	PP2068 : and2 port map (X(0), Y(39), N0_39_39);
	-- signal N0_39_40 : std_logic;
	PP2069 : and2 port map (X(1), Y(39), N0_39_40);
	-- signal N0_39_41 : std_logic;
	PP2070 : and2 port map (X(2), Y(39), N0_39_41);
	-- signal N0_39_42 : std_logic;
	PP2071 : and2 port map (X(3), Y(39), N0_39_42);
	-- signal N0_39_43 : std_logic;
	PP2072 : and2 port map (X(4), Y(39), N0_39_43);
	-- signal N0_39_44 : std_logic;
	PP2073 : and2 port map (X(5), Y(39), N0_39_44);
	-- signal N0_39_45 : std_logic;
	PP2074 : and2 port map (X(6), Y(39), N0_39_45);
	-- signal N0_39_46 : std_logic;
	PP2075 : and2 port map (X(7), Y(39), N0_39_46);
	-- signal N0_39_47 : std_logic;
	PP2076 : and2 port map (X(8), Y(39), N0_39_47);
	-- signal N0_39_48 : std_logic;
	PP2077 : and2 port map (X(9), Y(39), N0_39_48);
	-- signal N0_39_49 : std_logic;
	PP2078 : and2 port map (X(10), Y(39), N0_39_49);
	-- signal N0_39_50 : std_logic;
	PP2079 : and2 port map (X(11), Y(39), N0_39_50);
	-- signal N0_39_51 : std_logic;
	PP2080 : and2 port map (X(12), Y(39), N0_39_51);
	-- signal N0_39_52 : std_logic;
	PP2081 : and2 port map (X(13), Y(39), N0_39_52);
	-- signal N0_39_53 : std_logic;
	PP2082 : and2 port map (X(14), Y(39), N0_39_53);
	-- signal N0_39_54 : std_logic;
	PP2083 : and2 port map (X(15), Y(39), N0_39_54);
	-- signal N0_39_55 : std_logic;
	PP2084 : and2 port map (X(16), Y(39), N0_39_55);
	-- signal N0_39_56 : std_logic;
	PP2085 : and2 port map (X(17), Y(39), N0_39_56);
	-- signal N0_39_57 : std_logic;
	PP2086 : and2 port map (X(18), Y(39), N0_39_57);
	-- signal N0_39_58 : std_logic;
	PP2087 : and2 port map (X(19), Y(39), N0_39_58);
	-- signal N0_39_59 : std_logic;
	PP2088 : and2 port map (X(20), Y(39), N0_39_59);
	-- signal N0_39_60 : std_logic;
	PP2089 : and2 port map (X(21), Y(39), N0_39_60);
	-- signal N0_39_61 : std_logic;
	PP2090 : and2 port map (X(22), Y(39), N0_39_61);
	-- signal N0_39_62 : std_logic;
	PP2091 : and2 port map (X(23), Y(39), N0_39_62);
	-- signal N0_39_63 : std_logic;
	PP2092 : and2 port map (X(24), Y(39), N0_39_63);
	-- signal N0_39_64 : std_logic;
	PP2093 : and2 port map (X(25), Y(39), N0_39_64);
	-- signal N0_39_65 : std_logic;
	PP2094 : and2 port map (X(26), Y(39), N0_39_65);
	-- signal N0_39_66 : std_logic;
	PP2095 : and2 port map (X(27), Y(39), N0_39_66);
	-- signal N0_39_67 : std_logic;
	PP2096 : and2 port map (X(28), Y(39), N0_39_67);
	-- signal N0_39_68 : std_logic;
	PP2097 : and2 port map (X(29), Y(39), N0_39_68);
	-- signal N0_39_69 : std_logic;
	PP2098 : and2 port map (X(30), Y(39), N0_39_69);
	-- signal N0_39_70 : std_logic;
	PP2099 : and2 port map (X(31), Y(39), N0_39_70);
	-- signal N0_39_71 : std_logic;
	PP2100 : and2 port map (X(32), Y(39), N0_39_71);
	-- signal N0_39_72 : std_logic;
	PP2101 : and2 port map (X(33), Y(39), N0_39_72);
	-- signal N0_39_73 : std_logic;
	PP2102 : and2 port map (X(34), Y(39), N0_39_73);
	-- signal N0_39_74 : std_logic;
	PP2103 : and2 port map (X(35), Y(39), N0_39_74);
	-- signal N0_39_75 : std_logic;
	PP2104 : and2 port map (X(36), Y(39), N0_39_75);
	-- signal N0_39_76 : std_logic;
	PP2105 : and2 port map (X(37), Y(39), N0_39_76);
	-- signal N0_39_77 : std_logic;
	PP2106 : and2 port map (X(38), Y(39), N0_39_77);
	-- signal N0_39_78 : std_logic;
	PP2107 : and2 port map (X(39), Y(39), N0_39_78);
	-- signal N0_39_79 : std_logic;
	PP2108 : and2 port map (X(40), Y(39), N0_39_79);
	-- signal N0_39_80 : std_logic;
	PP2109 : and2 port map (X(41), Y(39), N0_39_80);
	-- signal N0_39_81 : std_logic;
	PP2110 : and2 port map (X(42), Y(39), N0_39_81);
	-- signal N0_39_82 : std_logic;
	PP2111 : and2 port map (X(43), Y(39), N0_39_82);
	-- signal N0_39_83 : std_logic;
	PP2112 : and2 port map (X(44), Y(39), N0_39_83);
	-- signal N0_39_84 : std_logic;
	PP2113 : and2 port map (X(45), Y(39), N0_39_84);
	-- signal N0_39_85 : std_logic;
	PP2114 : and2 port map (X(46), Y(39), N0_39_85);
	-- signal N0_39_86 : std_logic;
	PP2115 : and2 port map (X(47), Y(39), N0_39_86);
	-- signal N0_39_87 : std_logic;
	PP2116 : and2 port map (X(48), Y(39), N0_39_87);
	-- signal N0_39_88 : std_logic;
	PP2117 : and2 port map (X(49), Y(39), N0_39_88);
	-- signal N0_39_89 : std_logic;
	PP2118 : and2 port map (X(50), Y(39), N0_39_89);
	-- signal N0_39_90 : std_logic;
	PP2119 : and2 port map (X(51), Y(39), N0_39_90);
	-- signal N0_39_91 : std_logic;
	PP2120 : and2 port map ('1', Y(39), N0_39_91);
	-- signal N0_40_40 : std_logic;
	PP2121 : and2 port map (X(0), Y(40), N0_40_40);
	-- signal N0_40_41 : std_logic;
	PP2122 : and2 port map (X(1), Y(40), N0_40_41);
	-- signal N0_40_42 : std_logic;
	PP2123 : and2 port map (X(2), Y(40), N0_40_42);
	-- signal N0_40_43 : std_logic;
	PP2124 : and2 port map (X(3), Y(40), N0_40_43);
	-- signal N0_40_44 : std_logic;
	PP2125 : and2 port map (X(4), Y(40), N0_40_44);
	-- signal N0_40_45 : std_logic;
	PP2126 : and2 port map (X(5), Y(40), N0_40_45);
	-- signal N0_40_46 : std_logic;
	PP2127 : and2 port map (X(6), Y(40), N0_40_46);
	-- signal N0_40_47 : std_logic;
	PP2128 : and2 port map (X(7), Y(40), N0_40_47);
	-- signal N0_40_48 : std_logic;
	PP2129 : and2 port map (X(8), Y(40), N0_40_48);
	-- signal N0_40_49 : std_logic;
	PP2130 : and2 port map (X(9), Y(40), N0_40_49);
	-- signal N0_40_50 : std_logic;
	PP2131 : and2 port map (X(10), Y(40), N0_40_50);
	-- signal N0_40_51 : std_logic;
	PP2132 : and2 port map (X(11), Y(40), N0_40_51);
	-- signal N0_40_52 : std_logic;
	PP2133 : and2 port map (X(12), Y(40), N0_40_52);
	-- signal N0_40_53 : std_logic;
	PP2134 : and2 port map (X(13), Y(40), N0_40_53);
	-- signal N0_40_54 : std_logic;
	PP2135 : and2 port map (X(14), Y(40), N0_40_54);
	-- signal N0_40_55 : std_logic;
	PP2136 : and2 port map (X(15), Y(40), N0_40_55);
	-- signal N0_40_56 : std_logic;
	PP2137 : and2 port map (X(16), Y(40), N0_40_56);
	-- signal N0_40_57 : std_logic;
	PP2138 : and2 port map (X(17), Y(40), N0_40_57);
	-- signal N0_40_58 : std_logic;
	PP2139 : and2 port map (X(18), Y(40), N0_40_58);
	-- signal N0_40_59 : std_logic;
	PP2140 : and2 port map (X(19), Y(40), N0_40_59);
	-- signal N0_40_60 : std_logic;
	PP2141 : and2 port map (X(20), Y(40), N0_40_60);
	-- signal N0_40_61 : std_logic;
	PP2142 : and2 port map (X(21), Y(40), N0_40_61);
	-- signal N0_40_62 : std_logic;
	PP2143 : and2 port map (X(22), Y(40), N0_40_62);
	-- signal N0_40_63 : std_logic;
	PP2144 : and2 port map (X(23), Y(40), N0_40_63);
	-- signal N0_40_64 : std_logic;
	PP2145 : and2 port map (X(24), Y(40), N0_40_64);
	-- signal N0_40_65 : std_logic;
	PP2146 : and2 port map (X(25), Y(40), N0_40_65);
	-- signal N0_40_66 : std_logic;
	PP2147 : and2 port map (X(26), Y(40), N0_40_66);
	-- signal N0_40_67 : std_logic;
	PP2148 : and2 port map (X(27), Y(40), N0_40_67);
	-- signal N0_40_68 : std_logic;
	PP2149 : and2 port map (X(28), Y(40), N0_40_68);
	-- signal N0_40_69 : std_logic;
	PP2150 : and2 port map (X(29), Y(40), N0_40_69);
	-- signal N0_40_70 : std_logic;
	PP2151 : and2 port map (X(30), Y(40), N0_40_70);
	-- signal N0_40_71 : std_logic;
	PP2152 : and2 port map (X(31), Y(40), N0_40_71);
	-- signal N0_40_72 : std_logic;
	PP2153 : and2 port map (X(32), Y(40), N0_40_72);
	-- signal N0_40_73 : std_logic;
	PP2154 : and2 port map (X(33), Y(40), N0_40_73);
	-- signal N0_40_74 : std_logic;
	PP2155 : and2 port map (X(34), Y(40), N0_40_74);
	-- signal N0_40_75 : std_logic;
	PP2156 : and2 port map (X(35), Y(40), N0_40_75);
	-- signal N0_40_76 : std_logic;
	PP2157 : and2 port map (X(36), Y(40), N0_40_76);
	-- signal N0_40_77 : std_logic;
	PP2158 : and2 port map (X(37), Y(40), N0_40_77);
	-- signal N0_40_78 : std_logic;
	PP2159 : and2 port map (X(38), Y(40), N0_40_78);
	-- signal N0_40_79 : std_logic;
	PP2160 : and2 port map (X(39), Y(40), N0_40_79);
	-- signal N0_40_80 : std_logic;
	PP2161 : and2 port map (X(40), Y(40), N0_40_80);
	-- signal N0_40_81 : std_logic;
	PP2162 : and2 port map (X(41), Y(40), N0_40_81);
	-- signal N0_40_82 : std_logic;
	PP2163 : and2 port map (X(42), Y(40), N0_40_82);
	-- signal N0_40_83 : std_logic;
	PP2164 : and2 port map (X(43), Y(40), N0_40_83);
	-- signal N0_40_84 : std_logic;
	PP2165 : and2 port map (X(44), Y(40), N0_40_84);
	-- signal N0_40_85 : std_logic;
	PP2166 : and2 port map (X(45), Y(40), N0_40_85);
	-- signal N0_40_86 : std_logic;
	PP2167 : and2 port map (X(46), Y(40), N0_40_86);
	-- signal N0_40_87 : std_logic;
	PP2168 : and2 port map (X(47), Y(40), N0_40_87);
	-- signal N0_40_88 : std_logic;
	PP2169 : and2 port map (X(48), Y(40), N0_40_88);
	-- signal N0_40_89 : std_logic;
	PP2170 : and2 port map (X(49), Y(40), N0_40_89);
	-- signal N0_40_90 : std_logic;
	PP2171 : and2 port map (X(50), Y(40), N0_40_90);
	-- signal N0_40_91 : std_logic;
	PP2172 : and2 port map (X(51), Y(40), N0_40_91);
	-- signal N0_40_92 : std_logic;
	PP2173 : and2 port map ('1', Y(40), N0_40_92);
	-- signal N0_41_41 : std_logic;
	PP2174 : and2 port map (X(0), Y(41), N0_41_41);
	-- signal N0_41_42 : std_logic;
	PP2175 : and2 port map (X(1), Y(41), N0_41_42);
	-- signal N0_41_43 : std_logic;
	PP2176 : and2 port map (X(2), Y(41), N0_41_43);
	-- signal N0_41_44 : std_logic;
	PP2177 : and2 port map (X(3), Y(41), N0_41_44);
	-- signal N0_41_45 : std_logic;
	PP2178 : and2 port map (X(4), Y(41), N0_41_45);
	-- signal N0_41_46 : std_logic;
	PP2179 : and2 port map (X(5), Y(41), N0_41_46);
	-- signal N0_41_47 : std_logic;
	PP2180 : and2 port map (X(6), Y(41), N0_41_47);
	-- signal N0_41_48 : std_logic;
	PP2181 : and2 port map (X(7), Y(41), N0_41_48);
	-- signal N0_41_49 : std_logic;
	PP2182 : and2 port map (X(8), Y(41), N0_41_49);
	-- signal N0_41_50 : std_logic;
	PP2183 : and2 port map (X(9), Y(41), N0_41_50);
	-- signal N0_41_51 : std_logic;
	PP2184 : and2 port map (X(10), Y(41), N0_41_51);
	-- signal N0_41_52 : std_logic;
	PP2185 : and2 port map (X(11), Y(41), N0_41_52);
	-- signal N0_41_53 : std_logic;
	PP2186 : and2 port map (X(12), Y(41), N0_41_53);
	-- signal N0_41_54 : std_logic;
	PP2187 : and2 port map (X(13), Y(41), N0_41_54);
	-- signal N0_41_55 : std_logic;
	PP2188 : and2 port map (X(14), Y(41), N0_41_55);
	-- signal N0_41_56 : std_logic;
	PP2189 : and2 port map (X(15), Y(41), N0_41_56);
	-- signal N0_41_57 : std_logic;
	PP2190 : and2 port map (X(16), Y(41), N0_41_57);
	-- signal N0_41_58 : std_logic;
	PP2191 : and2 port map (X(17), Y(41), N0_41_58);
	-- signal N0_41_59 : std_logic;
	PP2192 : and2 port map (X(18), Y(41), N0_41_59);
	-- signal N0_41_60 : std_logic;
	PP2193 : and2 port map (X(19), Y(41), N0_41_60);
	-- signal N0_41_61 : std_logic;
	PP2194 : and2 port map (X(20), Y(41), N0_41_61);
	-- signal N0_41_62 : std_logic;
	PP2195 : and2 port map (X(21), Y(41), N0_41_62);
	-- signal N0_41_63 : std_logic;
	PP2196 : and2 port map (X(22), Y(41), N0_41_63);
	-- signal N0_41_64 : std_logic;
	PP2197 : and2 port map (X(23), Y(41), N0_41_64);
	-- signal N0_41_65 : std_logic;
	PP2198 : and2 port map (X(24), Y(41), N0_41_65);
	-- signal N0_41_66 : std_logic;
	PP2199 : and2 port map (X(25), Y(41), N0_41_66);
	-- signal N0_41_67 : std_logic;
	PP2200 : and2 port map (X(26), Y(41), N0_41_67);
	-- signal N0_41_68 : std_logic;
	PP2201 : and2 port map (X(27), Y(41), N0_41_68);
	-- signal N0_41_69 : std_logic;
	PP2202 : and2 port map (X(28), Y(41), N0_41_69);
	-- signal N0_41_70 : std_logic;
	PP2203 : and2 port map (X(29), Y(41), N0_41_70);
	-- signal N0_41_71 : std_logic;
	PP2204 : and2 port map (X(30), Y(41), N0_41_71);
	-- signal N0_41_72 : std_logic;
	PP2205 : and2 port map (X(31), Y(41), N0_41_72);
	-- signal N0_41_73 : std_logic;
	PP2206 : and2 port map (X(32), Y(41), N0_41_73);
	-- signal N0_41_74 : std_logic;
	PP2207 : and2 port map (X(33), Y(41), N0_41_74);
	-- signal N0_41_75 : std_logic;
	PP2208 : and2 port map (X(34), Y(41), N0_41_75);
	-- signal N0_41_76 : std_logic;
	PP2209 : and2 port map (X(35), Y(41), N0_41_76);
	-- signal N0_41_77 : std_logic;
	PP2210 : and2 port map (X(36), Y(41), N0_41_77);
	-- signal N0_41_78 : std_logic;
	PP2211 : and2 port map (X(37), Y(41), N0_41_78);
	-- signal N0_41_79 : std_logic;
	PP2212 : and2 port map (X(38), Y(41), N0_41_79);
	-- signal N0_41_80 : std_logic;
	PP2213 : and2 port map (X(39), Y(41), N0_41_80);
	-- signal N0_41_81 : std_logic;
	PP2214 : and2 port map (X(40), Y(41), N0_41_81);
	-- signal N0_41_82 : std_logic;
	PP2215 : and2 port map (X(41), Y(41), N0_41_82);
	-- signal N0_41_83 : std_logic;
	PP2216 : and2 port map (X(42), Y(41), N0_41_83);
	-- signal N0_41_84 : std_logic;
	PP2217 : and2 port map (X(43), Y(41), N0_41_84);
	-- signal N0_41_85 : std_logic;
	PP2218 : and2 port map (X(44), Y(41), N0_41_85);
	-- signal N0_41_86 : std_logic;
	PP2219 : and2 port map (X(45), Y(41), N0_41_86);
	-- signal N0_41_87 : std_logic;
	PP2220 : and2 port map (X(46), Y(41), N0_41_87);
	-- signal N0_41_88 : std_logic;
	PP2221 : and2 port map (X(47), Y(41), N0_41_88);
	-- signal N0_41_89 : std_logic;
	PP2222 : and2 port map (X(48), Y(41), N0_41_89);
	-- signal N0_41_90 : std_logic;
	PP2223 : and2 port map (X(49), Y(41), N0_41_90);
	-- signal N0_41_91 : std_logic;
	PP2224 : and2 port map (X(50), Y(41), N0_41_91);
	-- signal N0_41_92 : std_logic;
	PP2225 : and2 port map (X(51), Y(41), N0_41_92);
	-- signal N0_41_93 : std_logic;
	PP2226 : and2 port map ('1', Y(41), N0_41_93);
	-- signal N0_42_42 : std_logic;
	PP2227 : and2 port map (X(0), Y(42), N0_42_42);
	-- signal N0_42_43 : std_logic;
	PP2228 : and2 port map (X(1), Y(42), N0_42_43);
	-- signal N0_42_44 : std_logic;
	PP2229 : and2 port map (X(2), Y(42), N0_42_44);
	-- signal N0_42_45 : std_logic;
	PP2230 : and2 port map (X(3), Y(42), N0_42_45);
	-- signal N0_42_46 : std_logic;
	PP2231 : and2 port map (X(4), Y(42), N0_42_46);
	-- signal N0_42_47 : std_logic;
	PP2232 : and2 port map (X(5), Y(42), N0_42_47);
	-- signal N0_42_48 : std_logic;
	PP2233 : and2 port map (X(6), Y(42), N0_42_48);
	-- signal N0_42_49 : std_logic;
	PP2234 : and2 port map (X(7), Y(42), N0_42_49);
	-- signal N0_42_50 : std_logic;
	PP2235 : and2 port map (X(8), Y(42), N0_42_50);
	-- signal N0_42_51 : std_logic;
	PP2236 : and2 port map (X(9), Y(42), N0_42_51);
	-- signal N0_42_52 : std_logic;
	PP2237 : and2 port map (X(10), Y(42), N0_42_52);
	-- signal N0_42_53 : std_logic;
	PP2238 : and2 port map (X(11), Y(42), N0_42_53);
	-- signal N0_42_54 : std_logic;
	PP2239 : and2 port map (X(12), Y(42), N0_42_54);
	-- signal N0_42_55 : std_logic;
	PP2240 : and2 port map (X(13), Y(42), N0_42_55);
	-- signal N0_42_56 : std_logic;
	PP2241 : and2 port map (X(14), Y(42), N0_42_56);
	-- signal N0_42_57 : std_logic;
	PP2242 : and2 port map (X(15), Y(42), N0_42_57);
	-- signal N0_42_58 : std_logic;
	PP2243 : and2 port map (X(16), Y(42), N0_42_58);
	-- signal N0_42_59 : std_logic;
	PP2244 : and2 port map (X(17), Y(42), N0_42_59);
	-- signal N0_42_60 : std_logic;
	PP2245 : and2 port map (X(18), Y(42), N0_42_60);
	-- signal N0_42_61 : std_logic;
	PP2246 : and2 port map (X(19), Y(42), N0_42_61);
	-- signal N0_42_62 : std_logic;
	PP2247 : and2 port map (X(20), Y(42), N0_42_62);
	-- signal N0_42_63 : std_logic;
	PP2248 : and2 port map (X(21), Y(42), N0_42_63);
	-- signal N0_42_64 : std_logic;
	PP2249 : and2 port map (X(22), Y(42), N0_42_64);
	-- signal N0_42_65 : std_logic;
	PP2250 : and2 port map (X(23), Y(42), N0_42_65);
	-- signal N0_42_66 : std_logic;
	PP2251 : and2 port map (X(24), Y(42), N0_42_66);
	-- signal N0_42_67 : std_logic;
	PP2252 : and2 port map (X(25), Y(42), N0_42_67);
	-- signal N0_42_68 : std_logic;
	PP2253 : and2 port map (X(26), Y(42), N0_42_68);
	-- signal N0_42_69 : std_logic;
	PP2254 : and2 port map (X(27), Y(42), N0_42_69);
	-- signal N0_42_70 : std_logic;
	PP2255 : and2 port map (X(28), Y(42), N0_42_70);
	-- signal N0_42_71 : std_logic;
	PP2256 : and2 port map (X(29), Y(42), N0_42_71);
	-- signal N0_42_72 : std_logic;
	PP2257 : and2 port map (X(30), Y(42), N0_42_72);
	-- signal N0_42_73 : std_logic;
	PP2258 : and2 port map (X(31), Y(42), N0_42_73);
	-- signal N0_42_74 : std_logic;
	PP2259 : and2 port map (X(32), Y(42), N0_42_74);
	-- signal N0_42_75 : std_logic;
	PP2260 : and2 port map (X(33), Y(42), N0_42_75);
	-- signal N0_42_76 : std_logic;
	PP2261 : and2 port map (X(34), Y(42), N0_42_76);
	-- signal N0_42_77 : std_logic;
	PP2262 : and2 port map (X(35), Y(42), N0_42_77);
	-- signal N0_42_78 : std_logic;
	PP2263 : and2 port map (X(36), Y(42), N0_42_78);
	-- signal N0_42_79 : std_logic;
	PP2264 : and2 port map (X(37), Y(42), N0_42_79);
	-- signal N0_42_80 : std_logic;
	PP2265 : and2 port map (X(38), Y(42), N0_42_80);
	-- signal N0_42_81 : std_logic;
	PP2266 : and2 port map (X(39), Y(42), N0_42_81);
	-- signal N0_42_82 : std_logic;
	PP2267 : and2 port map (X(40), Y(42), N0_42_82);
	-- signal N0_42_83 : std_logic;
	PP2268 : and2 port map (X(41), Y(42), N0_42_83);
	-- signal N0_42_84 : std_logic;
	PP2269 : and2 port map (X(42), Y(42), N0_42_84);
	-- signal N0_42_85 : std_logic;
	PP2270 : and2 port map (X(43), Y(42), N0_42_85);
	-- signal N0_42_86 : std_logic;
	PP2271 : and2 port map (X(44), Y(42), N0_42_86);
	-- signal N0_42_87 : std_logic;
	PP2272 : and2 port map (X(45), Y(42), N0_42_87);
	-- signal N0_42_88 : std_logic;
	PP2273 : and2 port map (X(46), Y(42), N0_42_88);
	-- signal N0_42_89 : std_logic;
	PP2274 : and2 port map (X(47), Y(42), N0_42_89);
	-- signal N0_42_90 : std_logic;
	PP2275 : and2 port map (X(48), Y(42), N0_42_90);
	-- signal N0_42_91 : std_logic;
	PP2276 : and2 port map (X(49), Y(42), N0_42_91);
	-- signal N0_42_92 : std_logic;
	PP2277 : and2 port map (X(50), Y(42), N0_42_92);
	-- signal N0_42_93 : std_logic;
	PP2278 : and2 port map (X(51), Y(42), N0_42_93);
	-- signal N0_42_94 : std_logic;
	PP2279 : and2 port map ('1', Y(42), N0_42_94);
	-- signal N0_43_43 : std_logic;
	PP2280 : and2 port map (X(0), Y(43), N0_43_43);
	-- signal N0_43_44 : std_logic;
	PP2281 : and2 port map (X(1), Y(43), N0_43_44);
	-- signal N0_43_45 : std_logic;
	PP2282 : and2 port map (X(2), Y(43), N0_43_45);
	-- signal N0_43_46 : std_logic;
	PP2283 : and2 port map (X(3), Y(43), N0_43_46);
	-- signal N0_43_47 : std_logic;
	PP2284 : and2 port map (X(4), Y(43), N0_43_47);
	-- signal N0_43_48 : std_logic;
	PP2285 : and2 port map (X(5), Y(43), N0_43_48);
	-- signal N0_43_49 : std_logic;
	PP2286 : and2 port map (X(6), Y(43), N0_43_49);
	-- signal N0_43_50 : std_logic;
	PP2287 : and2 port map (X(7), Y(43), N0_43_50);
	-- signal N0_43_51 : std_logic;
	PP2288 : and2 port map (X(8), Y(43), N0_43_51);
	-- signal N0_43_52 : std_logic;
	PP2289 : and2 port map (X(9), Y(43), N0_43_52);
	-- signal N0_43_53 : std_logic;
	PP2290 : and2 port map (X(10), Y(43), N0_43_53);
	-- signal N0_43_54 : std_logic;
	PP2291 : and2 port map (X(11), Y(43), N0_43_54);
	-- signal N0_43_55 : std_logic;
	PP2292 : and2 port map (X(12), Y(43), N0_43_55);
	-- signal N0_43_56 : std_logic;
	PP2293 : and2 port map (X(13), Y(43), N0_43_56);
	-- signal N0_43_57 : std_logic;
	PP2294 : and2 port map (X(14), Y(43), N0_43_57);
	-- signal N0_43_58 : std_logic;
	PP2295 : and2 port map (X(15), Y(43), N0_43_58);
	-- signal N0_43_59 : std_logic;
	PP2296 : and2 port map (X(16), Y(43), N0_43_59);
	-- signal N0_43_60 : std_logic;
	PP2297 : and2 port map (X(17), Y(43), N0_43_60);
	-- signal N0_43_61 : std_logic;
	PP2298 : and2 port map (X(18), Y(43), N0_43_61);
	-- signal N0_43_62 : std_logic;
	PP2299 : and2 port map (X(19), Y(43), N0_43_62);
	-- signal N0_43_63 : std_logic;
	PP2300 : and2 port map (X(20), Y(43), N0_43_63);
	-- signal N0_43_64 : std_logic;
	PP2301 : and2 port map (X(21), Y(43), N0_43_64);
	-- signal N0_43_65 : std_logic;
	PP2302 : and2 port map (X(22), Y(43), N0_43_65);
	-- signal N0_43_66 : std_logic;
	PP2303 : and2 port map (X(23), Y(43), N0_43_66);
	-- signal N0_43_67 : std_logic;
	PP2304 : and2 port map (X(24), Y(43), N0_43_67);
	-- signal N0_43_68 : std_logic;
	PP2305 : and2 port map (X(25), Y(43), N0_43_68);
	-- signal N0_43_69 : std_logic;
	PP2306 : and2 port map (X(26), Y(43), N0_43_69);
	-- signal N0_43_70 : std_logic;
	PP2307 : and2 port map (X(27), Y(43), N0_43_70);
	-- signal N0_43_71 : std_logic;
	PP2308 : and2 port map (X(28), Y(43), N0_43_71);
	-- signal N0_43_72 : std_logic;
	PP2309 : and2 port map (X(29), Y(43), N0_43_72);
	-- signal N0_43_73 : std_logic;
	PP2310 : and2 port map (X(30), Y(43), N0_43_73);
	-- signal N0_43_74 : std_logic;
	PP2311 : and2 port map (X(31), Y(43), N0_43_74);
	-- signal N0_43_75 : std_logic;
	PP2312 : and2 port map (X(32), Y(43), N0_43_75);
	-- signal N0_43_76 : std_logic;
	PP2313 : and2 port map (X(33), Y(43), N0_43_76);
	-- signal N0_43_77 : std_logic;
	PP2314 : and2 port map (X(34), Y(43), N0_43_77);
	-- signal N0_43_78 : std_logic;
	PP2315 : and2 port map (X(35), Y(43), N0_43_78);
	-- signal N0_43_79 : std_logic;
	PP2316 : and2 port map (X(36), Y(43), N0_43_79);
	-- signal N0_43_80 : std_logic;
	PP2317 : and2 port map (X(37), Y(43), N0_43_80);
	-- signal N0_43_81 : std_logic;
	PP2318 : and2 port map (X(38), Y(43), N0_43_81);
	-- signal N0_43_82 : std_logic;
	PP2319 : and2 port map (X(39), Y(43), N0_43_82);
	-- signal N0_43_83 : std_logic;
	PP2320 : and2 port map (X(40), Y(43), N0_43_83);
	-- signal N0_43_84 : std_logic;
	PP2321 : and2 port map (X(41), Y(43), N0_43_84);
	-- signal N0_43_85 : std_logic;
	PP2322 : and2 port map (X(42), Y(43), N0_43_85);
	-- signal N0_43_86 : std_logic;
	PP2323 : and2 port map (X(43), Y(43), N0_43_86);
	-- signal N0_43_87 : std_logic;
	PP2324 : and2 port map (X(44), Y(43), N0_43_87);
	-- signal N0_43_88 : std_logic;
	PP2325 : and2 port map (X(45), Y(43), N0_43_88);
	-- signal N0_43_89 : std_logic;
	PP2326 : and2 port map (X(46), Y(43), N0_43_89);
	-- signal N0_43_90 : std_logic;
	PP2327 : and2 port map (X(47), Y(43), N0_43_90);
	-- signal N0_43_91 : std_logic;
	PP2328 : and2 port map (X(48), Y(43), N0_43_91);
	-- signal N0_43_92 : std_logic;
	PP2329 : and2 port map (X(49), Y(43), N0_43_92);
	-- signal N0_43_93 : std_logic;
	PP2330 : and2 port map (X(50), Y(43), N0_43_93);
	-- signal N0_43_94 : std_logic;
	PP2331 : and2 port map (X(51), Y(43), N0_43_94);
	-- signal N0_43_95 : std_logic;
	PP2332 : and2 port map ('1', Y(43), N0_43_95);
	-- signal N0_44_44 : std_logic;
	PP2333 : and2 port map (X(0), Y(44), N0_44_44);
	-- signal N0_44_45 : std_logic;
	PP2334 : and2 port map (X(1), Y(44), N0_44_45);
	-- signal N0_44_46 : std_logic;
	PP2335 : and2 port map (X(2), Y(44), N0_44_46);
	-- signal N0_44_47 : std_logic;
	PP2336 : and2 port map (X(3), Y(44), N0_44_47);
	-- signal N0_44_48 : std_logic;
	PP2337 : and2 port map (X(4), Y(44), N0_44_48);
	-- signal N0_44_49 : std_logic;
	PP2338 : and2 port map (X(5), Y(44), N0_44_49);
	-- signal N0_44_50 : std_logic;
	PP2339 : and2 port map (X(6), Y(44), N0_44_50);
	-- signal N0_44_51 : std_logic;
	PP2340 : and2 port map (X(7), Y(44), N0_44_51);
	-- signal N0_44_52 : std_logic;
	PP2341 : and2 port map (X(8), Y(44), N0_44_52);
	-- signal N0_44_53 : std_logic;
	PP2342 : and2 port map (X(9), Y(44), N0_44_53);
	-- signal N0_44_54 : std_logic;
	PP2343 : and2 port map (X(10), Y(44), N0_44_54);
	-- signal N0_44_55 : std_logic;
	PP2344 : and2 port map (X(11), Y(44), N0_44_55);
	-- signal N0_44_56 : std_logic;
	PP2345 : and2 port map (X(12), Y(44), N0_44_56);
	-- signal N0_44_57 : std_logic;
	PP2346 : and2 port map (X(13), Y(44), N0_44_57);
	-- signal N0_44_58 : std_logic;
	PP2347 : and2 port map (X(14), Y(44), N0_44_58);
	-- signal N0_44_59 : std_logic;
	PP2348 : and2 port map (X(15), Y(44), N0_44_59);
	-- signal N0_44_60 : std_logic;
	PP2349 : and2 port map (X(16), Y(44), N0_44_60);
	-- signal N0_44_61 : std_logic;
	PP2350 : and2 port map (X(17), Y(44), N0_44_61);
	-- signal N0_44_62 : std_logic;
	PP2351 : and2 port map (X(18), Y(44), N0_44_62);
	-- signal N0_44_63 : std_logic;
	PP2352 : and2 port map (X(19), Y(44), N0_44_63);
	-- signal N0_44_64 : std_logic;
	PP2353 : and2 port map (X(20), Y(44), N0_44_64);
	-- signal N0_44_65 : std_logic;
	PP2354 : and2 port map (X(21), Y(44), N0_44_65);
	-- signal N0_44_66 : std_logic;
	PP2355 : and2 port map (X(22), Y(44), N0_44_66);
	-- signal N0_44_67 : std_logic;
	PP2356 : and2 port map (X(23), Y(44), N0_44_67);
	-- signal N0_44_68 : std_logic;
	PP2357 : and2 port map (X(24), Y(44), N0_44_68);
	-- signal N0_44_69 : std_logic;
	PP2358 : and2 port map (X(25), Y(44), N0_44_69);
	-- signal N0_44_70 : std_logic;
	PP2359 : and2 port map (X(26), Y(44), N0_44_70);
	-- signal N0_44_71 : std_logic;
	PP2360 : and2 port map (X(27), Y(44), N0_44_71);
	-- signal N0_44_72 : std_logic;
	PP2361 : and2 port map (X(28), Y(44), N0_44_72);
	-- signal N0_44_73 : std_logic;
	PP2362 : and2 port map (X(29), Y(44), N0_44_73);
	-- signal N0_44_74 : std_logic;
	PP2363 : and2 port map (X(30), Y(44), N0_44_74);
	-- signal N0_44_75 : std_logic;
	PP2364 : and2 port map (X(31), Y(44), N0_44_75);
	-- signal N0_44_76 : std_logic;
	PP2365 : and2 port map (X(32), Y(44), N0_44_76);
	-- signal N0_44_77 : std_logic;
	PP2366 : and2 port map (X(33), Y(44), N0_44_77);
	-- signal N0_44_78 : std_logic;
	PP2367 : and2 port map (X(34), Y(44), N0_44_78);
	-- signal N0_44_79 : std_logic;
	PP2368 : and2 port map (X(35), Y(44), N0_44_79);
	-- signal N0_44_80 : std_logic;
	PP2369 : and2 port map (X(36), Y(44), N0_44_80);
	-- signal N0_44_81 : std_logic;
	PP2370 : and2 port map (X(37), Y(44), N0_44_81);
	-- signal N0_44_82 : std_logic;
	PP2371 : and2 port map (X(38), Y(44), N0_44_82);
	-- signal N0_44_83 : std_logic;
	PP2372 : and2 port map (X(39), Y(44), N0_44_83);
	-- signal N0_44_84 : std_logic;
	PP2373 : and2 port map (X(40), Y(44), N0_44_84);
	-- signal N0_44_85 : std_logic;
	PP2374 : and2 port map (X(41), Y(44), N0_44_85);
	-- signal N0_44_86 : std_logic;
	PP2375 : and2 port map (X(42), Y(44), N0_44_86);
	-- signal N0_44_87 : std_logic;
	PP2376 : and2 port map (X(43), Y(44), N0_44_87);
	-- signal N0_44_88 : std_logic;
	PP2377 : and2 port map (X(44), Y(44), N0_44_88);
	-- signal N0_44_89 : std_logic;
	PP2378 : and2 port map (X(45), Y(44), N0_44_89);
	-- signal N0_44_90 : std_logic;
	PP2379 : and2 port map (X(46), Y(44), N0_44_90);
	-- signal N0_44_91 : std_logic;
	PP2380 : and2 port map (X(47), Y(44), N0_44_91);
	-- signal N0_44_92 : std_logic;
	PP2381 : and2 port map (X(48), Y(44), N0_44_92);
	-- signal N0_44_93 : std_logic;
	PP2382 : and2 port map (X(49), Y(44), N0_44_93);
	-- signal N0_44_94 : std_logic;
	PP2383 : and2 port map (X(50), Y(44), N0_44_94);
	-- signal N0_44_95 : std_logic;
	PP2384 : and2 port map (X(51), Y(44), N0_44_95);
	-- signal N0_44_96 : std_logic;
	PP2385 : and2 port map ('1', Y(44), N0_44_96);
	-- signal N0_45_45 : std_logic;
	PP2386 : and2 port map (X(0), Y(45), N0_45_45);
	-- signal N0_45_46 : std_logic;
	PP2387 : and2 port map (X(1), Y(45), N0_45_46);
	-- signal N0_45_47 : std_logic;
	PP2388 : and2 port map (X(2), Y(45), N0_45_47);
	-- signal N0_45_48 : std_logic;
	PP2389 : and2 port map (X(3), Y(45), N0_45_48);
	-- signal N0_45_49 : std_logic;
	PP2390 : and2 port map (X(4), Y(45), N0_45_49);
	-- signal N0_45_50 : std_logic;
	PP2391 : and2 port map (X(5), Y(45), N0_45_50);
	-- signal N0_45_51 : std_logic;
	PP2392 : and2 port map (X(6), Y(45), N0_45_51);
	-- signal N0_45_52 : std_logic;
	PP2393 : and2 port map (X(7), Y(45), N0_45_52);
	-- signal N0_45_53 : std_logic;
	PP2394 : and2 port map (X(8), Y(45), N0_45_53);
	-- signal N0_45_54 : std_logic;
	PP2395 : and2 port map (X(9), Y(45), N0_45_54);
	-- signal N0_45_55 : std_logic;
	PP2396 : and2 port map (X(10), Y(45), N0_45_55);
	-- signal N0_45_56 : std_logic;
	PP2397 : and2 port map (X(11), Y(45), N0_45_56);
	-- signal N0_45_57 : std_logic;
	PP2398 : and2 port map (X(12), Y(45), N0_45_57);
	-- signal N0_45_58 : std_logic;
	PP2399 : and2 port map (X(13), Y(45), N0_45_58);
	-- signal N0_45_59 : std_logic;
	PP2400 : and2 port map (X(14), Y(45), N0_45_59);
	-- signal N0_45_60 : std_logic;
	PP2401 : and2 port map (X(15), Y(45), N0_45_60);
	-- signal N0_45_61 : std_logic;
	PP2402 : and2 port map (X(16), Y(45), N0_45_61);
	-- signal N0_45_62 : std_logic;
	PP2403 : and2 port map (X(17), Y(45), N0_45_62);
	-- signal N0_45_63 : std_logic;
	PP2404 : and2 port map (X(18), Y(45), N0_45_63);
	-- signal N0_45_64 : std_logic;
	PP2405 : and2 port map (X(19), Y(45), N0_45_64);
	-- signal N0_45_65 : std_logic;
	PP2406 : and2 port map (X(20), Y(45), N0_45_65);
	-- signal N0_45_66 : std_logic;
	PP2407 : and2 port map (X(21), Y(45), N0_45_66);
	-- signal N0_45_67 : std_logic;
	PP2408 : and2 port map (X(22), Y(45), N0_45_67);
	-- signal N0_45_68 : std_logic;
	PP2409 : and2 port map (X(23), Y(45), N0_45_68);
	-- signal N0_45_69 : std_logic;
	PP2410 : and2 port map (X(24), Y(45), N0_45_69);
	-- signal N0_45_70 : std_logic;
	PP2411 : and2 port map (X(25), Y(45), N0_45_70);
	-- signal N0_45_71 : std_logic;
	PP2412 : and2 port map (X(26), Y(45), N0_45_71);
	-- signal N0_45_72 : std_logic;
	PP2413 : and2 port map (X(27), Y(45), N0_45_72);
	-- signal N0_45_73 : std_logic;
	PP2414 : and2 port map (X(28), Y(45), N0_45_73);
	-- signal N0_45_74 : std_logic;
	PP2415 : and2 port map (X(29), Y(45), N0_45_74);
	-- signal N0_45_75 : std_logic;
	PP2416 : and2 port map (X(30), Y(45), N0_45_75);
	-- signal N0_45_76 : std_logic;
	PP2417 : and2 port map (X(31), Y(45), N0_45_76);
	-- signal N0_45_77 : std_logic;
	PP2418 : and2 port map (X(32), Y(45), N0_45_77);
	-- signal N0_45_78 : std_logic;
	PP2419 : and2 port map (X(33), Y(45), N0_45_78);
	-- signal N0_45_79 : std_logic;
	PP2420 : and2 port map (X(34), Y(45), N0_45_79);
	-- signal N0_45_80 : std_logic;
	PP2421 : and2 port map (X(35), Y(45), N0_45_80);
	-- signal N0_45_81 : std_logic;
	PP2422 : and2 port map (X(36), Y(45), N0_45_81);
	-- signal N0_45_82 : std_logic;
	PP2423 : and2 port map (X(37), Y(45), N0_45_82);
	-- signal N0_45_83 : std_logic;
	PP2424 : and2 port map (X(38), Y(45), N0_45_83);
	-- signal N0_45_84 : std_logic;
	PP2425 : and2 port map (X(39), Y(45), N0_45_84);
	-- signal N0_45_85 : std_logic;
	PP2426 : and2 port map (X(40), Y(45), N0_45_85);
	-- signal N0_45_86 : std_logic;
	PP2427 : and2 port map (X(41), Y(45), N0_45_86);
	-- signal N0_45_87 : std_logic;
	PP2428 : and2 port map (X(42), Y(45), N0_45_87);
	-- signal N0_45_88 : std_logic;
	PP2429 : and2 port map (X(43), Y(45), N0_45_88);
	-- signal N0_45_89 : std_logic;
	PP2430 : and2 port map (X(44), Y(45), N0_45_89);
	-- signal N0_45_90 : std_logic;
	PP2431 : and2 port map (X(45), Y(45), N0_45_90);
	-- signal N0_45_91 : std_logic;
	PP2432 : and2 port map (X(46), Y(45), N0_45_91);
	-- signal N0_45_92 : std_logic;
	PP2433 : and2 port map (X(47), Y(45), N0_45_92);
	-- signal N0_45_93 : std_logic;
	PP2434 : and2 port map (X(48), Y(45), N0_45_93);
	-- signal N0_45_94 : std_logic;
	PP2435 : and2 port map (X(49), Y(45), N0_45_94);
	-- signal N0_45_95 : std_logic;
	PP2436 : and2 port map (X(50), Y(45), N0_45_95);
	-- signal N0_45_96 : std_logic;
	PP2437 : and2 port map (X(51), Y(45), N0_45_96);
	-- signal N0_45_97 : std_logic;
	PP2438 : and2 port map ('1', Y(45), N0_45_97);
	-- signal N0_46_46 : std_logic;
	PP2439 : and2 port map (X(0), Y(46), N0_46_46);
	-- signal N0_46_47 : std_logic;
	PP2440 : and2 port map (X(1), Y(46), N0_46_47);
	-- signal N0_46_48 : std_logic;
	PP2441 : and2 port map (X(2), Y(46), N0_46_48);
	-- signal N0_46_49 : std_logic;
	PP2442 : and2 port map (X(3), Y(46), N0_46_49);
	-- signal N0_46_50 : std_logic;
	PP2443 : and2 port map (X(4), Y(46), N0_46_50);
	-- signal N0_46_51 : std_logic;
	PP2444 : and2 port map (X(5), Y(46), N0_46_51);
	-- signal N0_46_52 : std_logic;
	PP2445 : and2 port map (X(6), Y(46), N0_46_52);
	-- signal N0_46_53 : std_logic;
	PP2446 : and2 port map (X(7), Y(46), N0_46_53);
	-- signal N0_46_54 : std_logic;
	PP2447 : and2 port map (X(8), Y(46), N0_46_54);
	-- signal N0_46_55 : std_logic;
	PP2448 : and2 port map (X(9), Y(46), N0_46_55);
	-- signal N0_46_56 : std_logic;
	PP2449 : and2 port map (X(10), Y(46), N0_46_56);
	-- signal N0_46_57 : std_logic;
	PP2450 : and2 port map (X(11), Y(46), N0_46_57);
	-- signal N0_46_58 : std_logic;
	PP2451 : and2 port map (X(12), Y(46), N0_46_58);
	-- signal N0_46_59 : std_logic;
	PP2452 : and2 port map (X(13), Y(46), N0_46_59);
	-- signal N0_46_60 : std_logic;
	PP2453 : and2 port map (X(14), Y(46), N0_46_60);
	-- signal N0_46_61 : std_logic;
	PP2454 : and2 port map (X(15), Y(46), N0_46_61);
	-- signal N0_46_62 : std_logic;
	PP2455 : and2 port map (X(16), Y(46), N0_46_62);
	-- signal N0_46_63 : std_logic;
	PP2456 : and2 port map (X(17), Y(46), N0_46_63);
	-- signal N0_46_64 : std_logic;
	PP2457 : and2 port map (X(18), Y(46), N0_46_64);
	-- signal N0_46_65 : std_logic;
	PP2458 : and2 port map (X(19), Y(46), N0_46_65);
	-- signal N0_46_66 : std_logic;
	PP2459 : and2 port map (X(20), Y(46), N0_46_66);
	-- signal N0_46_67 : std_logic;
	PP2460 : and2 port map (X(21), Y(46), N0_46_67);
	-- signal N0_46_68 : std_logic;
	PP2461 : and2 port map (X(22), Y(46), N0_46_68);
	-- signal N0_46_69 : std_logic;
	PP2462 : and2 port map (X(23), Y(46), N0_46_69);
	-- signal N0_46_70 : std_logic;
	PP2463 : and2 port map (X(24), Y(46), N0_46_70);
	-- signal N0_46_71 : std_logic;
	PP2464 : and2 port map (X(25), Y(46), N0_46_71);
	-- signal N0_46_72 : std_logic;
	PP2465 : and2 port map (X(26), Y(46), N0_46_72);
	-- signal N0_46_73 : std_logic;
	PP2466 : and2 port map (X(27), Y(46), N0_46_73);
	-- signal N0_46_74 : std_logic;
	PP2467 : and2 port map (X(28), Y(46), N0_46_74);
	-- signal N0_46_75 : std_logic;
	PP2468 : and2 port map (X(29), Y(46), N0_46_75);
	-- signal N0_46_76 : std_logic;
	PP2469 : and2 port map (X(30), Y(46), N0_46_76);
	-- signal N0_46_77 : std_logic;
	PP2470 : and2 port map (X(31), Y(46), N0_46_77);
	-- signal N0_46_78 : std_logic;
	PP2471 : and2 port map (X(32), Y(46), N0_46_78);
	-- signal N0_46_79 : std_logic;
	PP2472 : and2 port map (X(33), Y(46), N0_46_79);
	-- signal N0_46_80 : std_logic;
	PP2473 : and2 port map (X(34), Y(46), N0_46_80);
	-- signal N0_46_81 : std_logic;
	PP2474 : and2 port map (X(35), Y(46), N0_46_81);
	-- signal N0_46_82 : std_logic;
	PP2475 : and2 port map (X(36), Y(46), N0_46_82);
	-- signal N0_46_83 : std_logic;
	PP2476 : and2 port map (X(37), Y(46), N0_46_83);
	-- signal N0_46_84 : std_logic;
	PP2477 : and2 port map (X(38), Y(46), N0_46_84);
	-- signal N0_46_85 : std_logic;
	PP2478 : and2 port map (X(39), Y(46), N0_46_85);
	-- signal N0_46_86 : std_logic;
	PP2479 : and2 port map (X(40), Y(46), N0_46_86);
	-- signal N0_46_87 : std_logic;
	PP2480 : and2 port map (X(41), Y(46), N0_46_87);
	-- signal N0_46_88 : std_logic;
	PP2481 : and2 port map (X(42), Y(46), N0_46_88);
	-- signal N0_46_89 : std_logic;
	PP2482 : and2 port map (X(43), Y(46), N0_46_89);
	-- signal N0_46_90 : std_logic;
	PP2483 : and2 port map (X(44), Y(46), N0_46_90);
	-- signal N0_46_91 : std_logic;
	PP2484 : and2 port map (X(45), Y(46), N0_46_91);
	-- signal N0_46_92 : std_logic;
	PP2485 : and2 port map (X(46), Y(46), N0_46_92);
	-- signal N0_46_93 : std_logic;
	PP2486 : and2 port map (X(47), Y(46), N0_46_93);
	-- signal N0_46_94 : std_logic;
	PP2487 : and2 port map (X(48), Y(46), N0_46_94);
	-- signal N0_46_95 : std_logic;
	PP2488 : and2 port map (X(49), Y(46), N0_46_95);
	-- signal N0_46_96 : std_logic;
	PP2489 : and2 port map (X(50), Y(46), N0_46_96);
	-- signal N0_46_97 : std_logic;
	PP2490 : and2 port map (X(51), Y(46), N0_46_97);
	-- signal N0_46_98 : std_logic;
	PP2491 : and2 port map ('1', Y(46), N0_46_98);
	-- signal N0_47_47 : std_logic;
	PP2492 : and2 port map (X(0), Y(47), N0_47_47);
	-- signal N0_47_48 : std_logic;
	PP2493 : and2 port map (X(1), Y(47), N0_47_48);
	-- signal N0_47_49 : std_logic;
	PP2494 : and2 port map (X(2), Y(47), N0_47_49);
	-- signal N0_47_50 : std_logic;
	PP2495 : and2 port map (X(3), Y(47), N0_47_50);
	-- signal N0_47_51 : std_logic;
	PP2496 : and2 port map (X(4), Y(47), N0_47_51);
	-- signal N0_47_52 : std_logic;
	PP2497 : and2 port map (X(5), Y(47), N0_47_52);
	-- signal N0_47_53 : std_logic;
	PP2498 : and2 port map (X(6), Y(47), N0_47_53);
	-- signal N0_47_54 : std_logic;
	PP2499 : and2 port map (X(7), Y(47), N0_47_54);
	-- signal N0_47_55 : std_logic;
	PP2500 : and2 port map (X(8), Y(47), N0_47_55);
	-- signal N0_47_56 : std_logic;
	PP2501 : and2 port map (X(9), Y(47), N0_47_56);
	-- signal N0_47_57 : std_logic;
	PP2502 : and2 port map (X(10), Y(47), N0_47_57);
	-- signal N0_47_58 : std_logic;
	PP2503 : and2 port map (X(11), Y(47), N0_47_58);
	-- signal N0_47_59 : std_logic;
	PP2504 : and2 port map (X(12), Y(47), N0_47_59);
	-- signal N0_47_60 : std_logic;
	PP2505 : and2 port map (X(13), Y(47), N0_47_60);
	-- signal N0_47_61 : std_logic;
	PP2506 : and2 port map (X(14), Y(47), N0_47_61);
	-- signal N0_47_62 : std_logic;
	PP2507 : and2 port map (X(15), Y(47), N0_47_62);
	-- signal N0_47_63 : std_logic;
	PP2508 : and2 port map (X(16), Y(47), N0_47_63);
	-- signal N0_47_64 : std_logic;
	PP2509 : and2 port map (X(17), Y(47), N0_47_64);
	-- signal N0_47_65 : std_logic;
	PP2510 : and2 port map (X(18), Y(47), N0_47_65);
	-- signal N0_47_66 : std_logic;
	PP2511 : and2 port map (X(19), Y(47), N0_47_66);
	-- signal N0_47_67 : std_logic;
	PP2512 : and2 port map (X(20), Y(47), N0_47_67);
	-- signal N0_47_68 : std_logic;
	PP2513 : and2 port map (X(21), Y(47), N0_47_68);
	-- signal N0_47_69 : std_logic;
	PP2514 : and2 port map (X(22), Y(47), N0_47_69);
	-- signal N0_47_70 : std_logic;
	PP2515 : and2 port map (X(23), Y(47), N0_47_70);
	-- signal N0_47_71 : std_logic;
	PP2516 : and2 port map (X(24), Y(47), N0_47_71);
	-- signal N0_47_72 : std_logic;
	PP2517 : and2 port map (X(25), Y(47), N0_47_72);
	-- signal N0_47_73 : std_logic;
	PP2518 : and2 port map (X(26), Y(47), N0_47_73);
	-- signal N0_47_74 : std_logic;
	PP2519 : and2 port map (X(27), Y(47), N0_47_74);
	-- signal N0_47_75 : std_logic;
	PP2520 : and2 port map (X(28), Y(47), N0_47_75);
	-- signal N0_47_76 : std_logic;
	PP2521 : and2 port map (X(29), Y(47), N0_47_76);
	-- signal N0_47_77 : std_logic;
	PP2522 : and2 port map (X(30), Y(47), N0_47_77);
	-- signal N0_47_78 : std_logic;
	PP2523 : and2 port map (X(31), Y(47), N0_47_78);
	-- signal N0_47_79 : std_logic;
	PP2524 : and2 port map (X(32), Y(47), N0_47_79);
	-- signal N0_47_80 : std_logic;
	PP2525 : and2 port map (X(33), Y(47), N0_47_80);
	-- signal N0_47_81 : std_logic;
	PP2526 : and2 port map (X(34), Y(47), N0_47_81);
	-- signal N0_47_82 : std_logic;
	PP2527 : and2 port map (X(35), Y(47), N0_47_82);
	-- signal N0_47_83 : std_logic;
	PP2528 : and2 port map (X(36), Y(47), N0_47_83);
	-- signal N0_47_84 : std_logic;
	PP2529 : and2 port map (X(37), Y(47), N0_47_84);
	-- signal N0_47_85 : std_logic;
	PP2530 : and2 port map (X(38), Y(47), N0_47_85);
	-- signal N0_47_86 : std_logic;
	PP2531 : and2 port map (X(39), Y(47), N0_47_86);
	-- signal N0_47_87 : std_logic;
	PP2532 : and2 port map (X(40), Y(47), N0_47_87);
	-- signal N0_47_88 : std_logic;
	PP2533 : and2 port map (X(41), Y(47), N0_47_88);
	-- signal N0_47_89 : std_logic;
	PP2534 : and2 port map (X(42), Y(47), N0_47_89);
	-- signal N0_47_90 : std_logic;
	PP2535 : and2 port map (X(43), Y(47), N0_47_90);
	-- signal N0_47_91 : std_logic;
	PP2536 : and2 port map (X(44), Y(47), N0_47_91);
	-- signal N0_47_92 : std_logic;
	PP2537 : and2 port map (X(45), Y(47), N0_47_92);
	-- signal N0_47_93 : std_logic;
	PP2538 : and2 port map (X(46), Y(47), N0_47_93);
	-- signal N0_47_94 : std_logic;
	PP2539 : and2 port map (X(47), Y(47), N0_47_94);
	-- signal N0_47_95 : std_logic;
	PP2540 : and2 port map (X(48), Y(47), N0_47_95);
	-- signal N0_47_96 : std_logic;
	PP2541 : and2 port map (X(49), Y(47), N0_47_96);
	-- signal N0_47_97 : std_logic;
	PP2542 : and2 port map (X(50), Y(47), N0_47_97);
	-- signal N0_47_98 : std_logic;
	PP2543 : and2 port map (X(51), Y(47), N0_47_98);
	-- signal N0_47_99 : std_logic;
	PP2544 : and2 port map ('1', Y(47), N0_47_99);
	-- signal N0_48_48 : std_logic;
	PP2545 : and2 port map (X(0), Y(48), N0_48_48);
	-- signal N0_48_49 : std_logic;
	PP2546 : and2 port map (X(1), Y(48), N0_48_49);
	-- signal N0_48_50 : std_logic;
	PP2547 : and2 port map (X(2), Y(48), N0_48_50);
	-- signal N0_48_51 : std_logic;
	PP2548 : and2 port map (X(3), Y(48), N0_48_51);
	-- signal N0_48_52 : std_logic;
	PP2549 : and2 port map (X(4), Y(48), N0_48_52);
	-- signal N0_48_53 : std_logic;
	PP2550 : and2 port map (X(5), Y(48), N0_48_53);
	-- signal N0_48_54 : std_logic;
	PP2551 : and2 port map (X(6), Y(48), N0_48_54);
	-- signal N0_48_55 : std_logic;
	PP2552 : and2 port map (X(7), Y(48), N0_48_55);
	-- signal N0_48_56 : std_logic;
	PP2553 : and2 port map (X(8), Y(48), N0_48_56);
	-- signal N0_48_57 : std_logic;
	PP2554 : and2 port map (X(9), Y(48), N0_48_57);
	-- signal N0_48_58 : std_logic;
	PP2555 : and2 port map (X(10), Y(48), N0_48_58);
	-- signal N0_48_59 : std_logic;
	PP2556 : and2 port map (X(11), Y(48), N0_48_59);
	-- signal N0_48_60 : std_logic;
	PP2557 : and2 port map (X(12), Y(48), N0_48_60);
	-- signal N0_48_61 : std_logic;
	PP2558 : and2 port map (X(13), Y(48), N0_48_61);
	-- signal N0_48_62 : std_logic;
	PP2559 : and2 port map (X(14), Y(48), N0_48_62);
	-- signal N0_48_63 : std_logic;
	PP2560 : and2 port map (X(15), Y(48), N0_48_63);
	-- signal N0_48_64 : std_logic;
	PP2561 : and2 port map (X(16), Y(48), N0_48_64);
	-- signal N0_48_65 : std_logic;
	PP2562 : and2 port map (X(17), Y(48), N0_48_65);
	-- signal N0_48_66 : std_logic;
	PP2563 : and2 port map (X(18), Y(48), N0_48_66);
	-- signal N0_48_67 : std_logic;
	PP2564 : and2 port map (X(19), Y(48), N0_48_67);
	-- signal N0_48_68 : std_logic;
	PP2565 : and2 port map (X(20), Y(48), N0_48_68);
	-- signal N0_48_69 : std_logic;
	PP2566 : and2 port map (X(21), Y(48), N0_48_69);
	-- signal N0_48_70 : std_logic;
	PP2567 : and2 port map (X(22), Y(48), N0_48_70);
	-- signal N0_48_71 : std_logic;
	PP2568 : and2 port map (X(23), Y(48), N0_48_71);
	-- signal N0_48_72 : std_logic;
	PP2569 : and2 port map (X(24), Y(48), N0_48_72);
	-- signal N0_48_73 : std_logic;
	PP2570 : and2 port map (X(25), Y(48), N0_48_73);
	-- signal N0_48_74 : std_logic;
	PP2571 : and2 port map (X(26), Y(48), N0_48_74);
	-- signal N0_48_75 : std_logic;
	PP2572 : and2 port map (X(27), Y(48), N0_48_75);
	-- signal N0_48_76 : std_logic;
	PP2573 : and2 port map (X(28), Y(48), N0_48_76);
	-- signal N0_48_77 : std_logic;
	PP2574 : and2 port map (X(29), Y(48), N0_48_77);
	-- signal N0_48_78 : std_logic;
	PP2575 : and2 port map (X(30), Y(48), N0_48_78);
	-- signal N0_48_79 : std_logic;
	PP2576 : and2 port map (X(31), Y(48), N0_48_79);
	-- signal N0_48_80 : std_logic;
	PP2577 : and2 port map (X(32), Y(48), N0_48_80);
	-- signal N0_48_81 : std_logic;
	PP2578 : and2 port map (X(33), Y(48), N0_48_81);
	-- signal N0_48_82 : std_logic;
	PP2579 : and2 port map (X(34), Y(48), N0_48_82);
	-- signal N0_48_83 : std_logic;
	PP2580 : and2 port map (X(35), Y(48), N0_48_83);
	-- signal N0_48_84 : std_logic;
	PP2581 : and2 port map (X(36), Y(48), N0_48_84);
	-- signal N0_48_85 : std_logic;
	PP2582 : and2 port map (X(37), Y(48), N0_48_85);
	-- signal N0_48_86 : std_logic;
	PP2583 : and2 port map (X(38), Y(48), N0_48_86);
	-- signal N0_48_87 : std_logic;
	PP2584 : and2 port map (X(39), Y(48), N0_48_87);
	-- signal N0_48_88 : std_logic;
	PP2585 : and2 port map (X(40), Y(48), N0_48_88);
	-- signal N0_48_89 : std_logic;
	PP2586 : and2 port map (X(41), Y(48), N0_48_89);
	-- signal N0_48_90 : std_logic;
	PP2587 : and2 port map (X(42), Y(48), N0_48_90);
	-- signal N0_48_91 : std_logic;
	PP2588 : and2 port map (X(43), Y(48), N0_48_91);
	-- signal N0_48_92 : std_logic;
	PP2589 : and2 port map (X(44), Y(48), N0_48_92);
	-- signal N0_48_93 : std_logic;
	PP2590 : and2 port map (X(45), Y(48), N0_48_93);
	-- signal N0_48_94 : std_logic;
	PP2591 : and2 port map (X(46), Y(48), N0_48_94);
	-- signal N0_48_95 : std_logic;
	PP2592 : and2 port map (X(47), Y(48), N0_48_95);
	-- signal N0_48_96 : std_logic;
	PP2593 : and2 port map (X(48), Y(48), N0_48_96);
	-- signal N0_48_97 : std_logic;
	PP2594 : and2 port map (X(49), Y(48), N0_48_97);
	-- signal N0_48_98 : std_logic;
	PP2595 : and2 port map (X(50), Y(48), N0_48_98);
	-- signal N0_48_99 : std_logic;
	PP2596 : and2 port map (X(51), Y(48), N0_48_99);
	-- signal N0_48_100 : std_logic;
	PP2597 : and2 port map ('1', Y(48), N0_48_100);
	-- signal N0_49_49 : std_logic;
	PP2598 : and2 port map (X(0), Y(49), N0_49_49);
	-- signal N0_49_50 : std_logic;
	PP2599 : and2 port map (X(1), Y(49), N0_49_50);
	-- signal N0_49_51 : std_logic;
	PP2600 : and2 port map (X(2), Y(49), N0_49_51);
	-- signal N0_49_52 : std_logic;
	PP2601 : and2 port map (X(3), Y(49), N0_49_52);
	-- signal N0_49_53 : std_logic;
	PP2602 : and2 port map (X(4), Y(49), N0_49_53);
	-- signal N0_49_54 : std_logic;
	PP2603 : and2 port map (X(5), Y(49), N0_49_54);
	-- signal N0_49_55 : std_logic;
	PP2604 : and2 port map (X(6), Y(49), N0_49_55);
	-- signal N0_49_56 : std_logic;
	PP2605 : and2 port map (X(7), Y(49), N0_49_56);
	-- signal N0_49_57 : std_logic;
	PP2606 : and2 port map (X(8), Y(49), N0_49_57);
	-- signal N0_49_58 : std_logic;
	PP2607 : and2 port map (X(9), Y(49), N0_49_58);
	-- signal N0_49_59 : std_logic;
	PP2608 : and2 port map (X(10), Y(49), N0_49_59);
	-- signal N0_49_60 : std_logic;
	PP2609 : and2 port map (X(11), Y(49), N0_49_60);
	-- signal N0_49_61 : std_logic;
	PP2610 : and2 port map (X(12), Y(49), N0_49_61);
	-- signal N0_49_62 : std_logic;
	PP2611 : and2 port map (X(13), Y(49), N0_49_62);
	-- signal N0_49_63 : std_logic;
	PP2612 : and2 port map (X(14), Y(49), N0_49_63);
	-- signal N0_49_64 : std_logic;
	PP2613 : and2 port map (X(15), Y(49), N0_49_64);
	-- signal N0_49_65 : std_logic;
	PP2614 : and2 port map (X(16), Y(49), N0_49_65);
	-- signal N0_49_66 : std_logic;
	PP2615 : and2 port map (X(17), Y(49), N0_49_66);
	-- signal N0_49_67 : std_logic;
	PP2616 : and2 port map (X(18), Y(49), N0_49_67);
	-- signal N0_49_68 : std_logic;
	PP2617 : and2 port map (X(19), Y(49), N0_49_68);
	-- signal N0_49_69 : std_logic;
	PP2618 : and2 port map (X(20), Y(49), N0_49_69);
	-- signal N0_49_70 : std_logic;
	PP2619 : and2 port map (X(21), Y(49), N0_49_70);
	-- signal N0_49_71 : std_logic;
	PP2620 : and2 port map (X(22), Y(49), N0_49_71);
	-- signal N0_49_72 : std_logic;
	PP2621 : and2 port map (X(23), Y(49), N0_49_72);
	-- signal N0_49_73 : std_logic;
	PP2622 : and2 port map (X(24), Y(49), N0_49_73);
	-- signal N0_49_74 : std_logic;
	PP2623 : and2 port map (X(25), Y(49), N0_49_74);
	-- signal N0_49_75 : std_logic;
	PP2624 : and2 port map (X(26), Y(49), N0_49_75);
	-- signal N0_49_76 : std_logic;
	PP2625 : and2 port map (X(27), Y(49), N0_49_76);
	-- signal N0_49_77 : std_logic;
	PP2626 : and2 port map (X(28), Y(49), N0_49_77);
	-- signal N0_49_78 : std_logic;
	PP2627 : and2 port map (X(29), Y(49), N0_49_78);
	-- signal N0_49_79 : std_logic;
	PP2628 : and2 port map (X(30), Y(49), N0_49_79);
	-- signal N0_49_80 : std_logic;
	PP2629 : and2 port map (X(31), Y(49), N0_49_80);
	-- signal N0_49_81 : std_logic;
	PP2630 : and2 port map (X(32), Y(49), N0_49_81);
	-- signal N0_49_82 : std_logic;
	PP2631 : and2 port map (X(33), Y(49), N0_49_82);
	-- signal N0_49_83 : std_logic;
	PP2632 : and2 port map (X(34), Y(49), N0_49_83);
	-- signal N0_49_84 : std_logic;
	PP2633 : and2 port map (X(35), Y(49), N0_49_84);
	-- signal N0_49_85 : std_logic;
	PP2634 : and2 port map (X(36), Y(49), N0_49_85);
	-- signal N0_49_86 : std_logic;
	PP2635 : and2 port map (X(37), Y(49), N0_49_86);
	-- signal N0_49_87 : std_logic;
	PP2636 : and2 port map (X(38), Y(49), N0_49_87);
	-- signal N0_49_88 : std_logic;
	PP2637 : and2 port map (X(39), Y(49), N0_49_88);
	-- signal N0_49_89 : std_logic;
	PP2638 : and2 port map (X(40), Y(49), N0_49_89);
	-- signal N0_49_90 : std_logic;
	PP2639 : and2 port map (X(41), Y(49), N0_49_90);
	-- signal N0_49_91 : std_logic;
	PP2640 : and2 port map (X(42), Y(49), N0_49_91);
	-- signal N0_49_92 : std_logic;
	PP2641 : and2 port map (X(43), Y(49), N0_49_92);
	-- signal N0_49_93 : std_logic;
	PP2642 : and2 port map (X(44), Y(49), N0_49_93);
	-- signal N0_49_94 : std_logic;
	PP2643 : and2 port map (X(45), Y(49), N0_49_94);
	-- signal N0_49_95 : std_logic;
	PP2644 : and2 port map (X(46), Y(49), N0_49_95);
	-- signal N0_49_96 : std_logic;
	PP2645 : and2 port map (X(47), Y(49), N0_49_96);
	-- signal N0_49_97 : std_logic;
	PP2646 : and2 port map (X(48), Y(49), N0_49_97);
	-- signal N0_49_98 : std_logic;
	PP2647 : and2 port map (X(49), Y(49), N0_49_98);
	-- signal N0_49_99 : std_logic;
	PP2648 : and2 port map (X(50), Y(49), N0_49_99);
	-- signal N0_49_100 : std_logic;
	PP2649 : and2 port map (X(51), Y(49), N0_49_100);
	-- signal N0_49_101 : std_logic;
	PP2650 : and2 port map ('1', Y(49), N0_49_101);
	-- signal N0_50_50 : std_logic;
	PP2651 : and2 port map (X(0), Y(50), N0_50_50);
	-- signal N0_50_51 : std_logic;
	PP2652 : and2 port map (X(1), Y(50), N0_50_51);
	-- signal N0_50_52 : std_logic;
	PP2653 : and2 port map (X(2), Y(50), N0_50_52);
	-- signal N0_50_53 : std_logic;
	PP2654 : and2 port map (X(3), Y(50), N0_50_53);
	-- signal N0_50_54 : std_logic;
	PP2655 : and2 port map (X(4), Y(50), N0_50_54);
	-- signal N0_50_55 : std_logic;
	PP2656 : and2 port map (X(5), Y(50), N0_50_55);
	-- signal N0_50_56 : std_logic;
	PP2657 : and2 port map (X(6), Y(50), N0_50_56);
	-- signal N0_50_57 : std_logic;
	PP2658 : and2 port map (X(7), Y(50), N0_50_57);
	-- signal N0_50_58 : std_logic;
	PP2659 : and2 port map (X(8), Y(50), N0_50_58);
	-- signal N0_50_59 : std_logic;
	PP2660 : and2 port map (X(9), Y(50), N0_50_59);
	-- signal N0_50_60 : std_logic;
	PP2661 : and2 port map (X(10), Y(50), N0_50_60);
	-- signal N0_50_61 : std_logic;
	PP2662 : and2 port map (X(11), Y(50), N0_50_61);
	-- signal N0_50_62 : std_logic;
	PP2663 : and2 port map (X(12), Y(50), N0_50_62);
	-- signal N0_50_63 : std_logic;
	PP2664 : and2 port map (X(13), Y(50), N0_50_63);
	-- signal N0_50_64 : std_logic;
	PP2665 : and2 port map (X(14), Y(50), N0_50_64);
	-- signal N0_50_65 : std_logic;
	PP2666 : and2 port map (X(15), Y(50), N0_50_65);
	-- signal N0_50_66 : std_logic;
	PP2667 : and2 port map (X(16), Y(50), N0_50_66);
	-- signal N0_50_67 : std_logic;
	PP2668 : and2 port map (X(17), Y(50), N0_50_67);
	-- signal N0_50_68 : std_logic;
	PP2669 : and2 port map (X(18), Y(50), N0_50_68);
	-- signal N0_50_69 : std_logic;
	PP2670 : and2 port map (X(19), Y(50), N0_50_69);
	-- signal N0_50_70 : std_logic;
	PP2671 : and2 port map (X(20), Y(50), N0_50_70);
	-- signal N0_50_71 : std_logic;
	PP2672 : and2 port map (X(21), Y(50), N0_50_71);
	-- signal N0_50_72 : std_logic;
	PP2673 : and2 port map (X(22), Y(50), N0_50_72);
	-- signal N0_50_73 : std_logic;
	PP2674 : and2 port map (X(23), Y(50), N0_50_73);
	-- signal N0_50_74 : std_logic;
	PP2675 : and2 port map (X(24), Y(50), N0_50_74);
	-- signal N0_50_75 : std_logic;
	PP2676 : and2 port map (X(25), Y(50), N0_50_75);
	-- signal N0_50_76 : std_logic;
	PP2677 : and2 port map (X(26), Y(50), N0_50_76);
	-- signal N0_50_77 : std_logic;
	PP2678 : and2 port map (X(27), Y(50), N0_50_77);
	-- signal N0_50_78 : std_logic;
	PP2679 : and2 port map (X(28), Y(50), N0_50_78);
	-- signal N0_50_79 : std_logic;
	PP2680 : and2 port map (X(29), Y(50), N0_50_79);
	-- signal N0_50_80 : std_logic;
	PP2681 : and2 port map (X(30), Y(50), N0_50_80);
	-- signal N0_50_81 : std_logic;
	PP2682 : and2 port map (X(31), Y(50), N0_50_81);
	-- signal N0_50_82 : std_logic;
	PP2683 : and2 port map (X(32), Y(50), N0_50_82);
	-- signal N0_50_83 : std_logic;
	PP2684 : and2 port map (X(33), Y(50), N0_50_83);
	-- signal N0_50_84 : std_logic;
	PP2685 : and2 port map (X(34), Y(50), N0_50_84);
	-- signal N0_50_85 : std_logic;
	PP2686 : and2 port map (X(35), Y(50), N0_50_85);
	-- signal N0_50_86 : std_logic;
	PP2687 : and2 port map (X(36), Y(50), N0_50_86);
	-- signal N0_50_87 : std_logic;
	PP2688 : and2 port map (X(37), Y(50), N0_50_87);
	-- signal N0_50_88 : std_logic;
	PP2689 : and2 port map (X(38), Y(50), N0_50_88);
	-- signal N0_50_89 : std_logic;
	PP2690 : and2 port map (X(39), Y(50), N0_50_89);
	-- signal N0_50_90 : std_logic;
	PP2691 : and2 port map (X(40), Y(50), N0_50_90);
	-- signal N0_50_91 : std_logic;
	PP2692 : and2 port map (X(41), Y(50), N0_50_91);
	-- signal N0_50_92 : std_logic;
	PP2693 : and2 port map (X(42), Y(50), N0_50_92);
	-- signal N0_50_93 : std_logic;
	PP2694 : and2 port map (X(43), Y(50), N0_50_93);
	-- signal N0_50_94 : std_logic;
	PP2695 : and2 port map (X(44), Y(50), N0_50_94);
	-- signal N0_50_95 : std_logic;
	PP2696 : and2 port map (X(45), Y(50), N0_50_95);
	-- signal N0_50_96 : std_logic;
	PP2697 : and2 port map (X(46), Y(50), N0_50_96);
	-- signal N0_50_97 : std_logic;
	PP2698 : and2 port map (X(47), Y(50), N0_50_97);
	-- signal N0_50_98 : std_logic;
	PP2699 : and2 port map (X(48), Y(50), N0_50_98);
	-- signal N0_50_99 : std_logic;
	PP2700 : and2 port map (X(49), Y(50), N0_50_99);
	-- signal N0_50_100 : std_logic;
	PP2701 : and2 port map (X(50), Y(50), N0_50_100);
	-- signal N0_50_101 : std_logic;
	PP2702 : and2 port map (X(51), Y(50), N0_50_101);
	-- signal N0_50_102 : std_logic;
	PP2703 : and2 port map ('1', Y(50), N0_50_102);
	-- signal N0_51_51 : std_logic;
	PP2704 : and2 port map (X(0), Y(51), N0_51_51);
	-- signal N0_51_52 : std_logic;
	PP2705 : and2 port map (X(1), Y(51), N0_51_52);
	-- signal N0_51_53 : std_logic;
	PP2706 : and2 port map (X(2), Y(51), N0_51_53);
	-- signal N0_51_54 : std_logic;
	PP2707 : and2 port map (X(3), Y(51), N0_51_54);
	-- signal N0_51_55 : std_logic;
	PP2708 : and2 port map (X(4), Y(51), N0_51_55);
	-- signal N0_51_56 : std_logic;
	PP2709 : and2 port map (X(5), Y(51), N0_51_56);
	-- signal N0_51_57 : std_logic;
	PP2710 : and2 port map (X(6), Y(51), N0_51_57);
	-- signal N0_51_58 : std_logic;
	PP2711 : and2 port map (X(7), Y(51), N0_51_58);
	-- signal N0_51_59 : std_logic;
	PP2712 : and2 port map (X(8), Y(51), N0_51_59);
	-- signal N0_51_60 : std_logic;
	PP2713 : and2 port map (X(9), Y(51), N0_51_60);
	-- signal N0_51_61 : std_logic;
	PP2714 : and2 port map (X(10), Y(51), N0_51_61);
	-- signal N0_51_62 : std_logic;
	PP2715 : and2 port map (X(11), Y(51), N0_51_62);
	-- signal N0_51_63 : std_logic;
	PP2716 : and2 port map (X(12), Y(51), N0_51_63);
	-- signal N0_51_64 : std_logic;
	PP2717 : and2 port map (X(13), Y(51), N0_51_64);
	-- signal N0_51_65 : std_logic;
	PP2718 : and2 port map (X(14), Y(51), N0_51_65);
	-- signal N0_51_66 : std_logic;
	PP2719 : and2 port map (X(15), Y(51), N0_51_66);
	-- signal N0_51_67 : std_logic;
	PP2720 : and2 port map (X(16), Y(51), N0_51_67);
	-- signal N0_51_68 : std_logic;
	PP2721 : and2 port map (X(17), Y(51), N0_51_68);
	-- signal N0_51_69 : std_logic;
	PP2722 : and2 port map (X(18), Y(51), N0_51_69);
	-- signal N0_51_70 : std_logic;
	PP2723 : and2 port map (X(19), Y(51), N0_51_70);
	-- signal N0_51_71 : std_logic;
	PP2724 : and2 port map (X(20), Y(51), N0_51_71);
	-- signal N0_51_72 : std_logic;
	PP2725 : and2 port map (X(21), Y(51), N0_51_72);
	-- signal N0_51_73 : std_logic;
	PP2726 : and2 port map (X(22), Y(51), N0_51_73);
	-- signal N0_51_74 : std_logic;
	PP2727 : and2 port map (X(23), Y(51), N0_51_74);
	-- signal N0_51_75 : std_logic;
	PP2728 : and2 port map (X(24), Y(51), N0_51_75);
	-- signal N0_51_76 : std_logic;
	PP2729 : and2 port map (X(25), Y(51), N0_51_76);
	-- signal N0_51_77 : std_logic;
	PP2730 : and2 port map (X(26), Y(51), N0_51_77);
	-- signal N0_51_78 : std_logic;
	PP2731 : and2 port map (X(27), Y(51), N0_51_78);
	-- signal N0_51_79 : std_logic;
	PP2732 : and2 port map (X(28), Y(51), N0_51_79);
	-- signal N0_51_80 : std_logic;
	PP2733 : and2 port map (X(29), Y(51), N0_51_80);
	-- signal N0_51_81 : std_logic;
	PP2734 : and2 port map (X(30), Y(51), N0_51_81);
	-- signal N0_51_82 : std_logic;
	PP2735 : and2 port map (X(31), Y(51), N0_51_82);
	-- signal N0_51_83 : std_logic;
	PP2736 : and2 port map (X(32), Y(51), N0_51_83);
	-- signal N0_51_84 : std_logic;
	PP2737 : and2 port map (X(33), Y(51), N0_51_84);
	-- signal N0_51_85 : std_logic;
	PP2738 : and2 port map (X(34), Y(51), N0_51_85);
	-- signal N0_51_86 : std_logic;
	PP2739 : and2 port map (X(35), Y(51), N0_51_86);
	-- signal N0_51_87 : std_logic;
	PP2740 : and2 port map (X(36), Y(51), N0_51_87);
	-- signal N0_51_88 : std_logic;
	PP2741 : and2 port map (X(37), Y(51), N0_51_88);
	-- signal N0_51_89 : std_logic;
	PP2742 : and2 port map (X(38), Y(51), N0_51_89);
	-- signal N0_51_90 : std_logic;
	PP2743 : and2 port map (X(39), Y(51), N0_51_90);
	-- signal N0_51_91 : std_logic;
	PP2744 : and2 port map (X(40), Y(51), N0_51_91);
	-- signal N0_51_92 : std_logic;
	PP2745 : and2 port map (X(41), Y(51), N0_51_92);
	-- signal N0_51_93 : std_logic;
	PP2746 : and2 port map (X(42), Y(51), N0_51_93);
	-- signal N0_51_94 : std_logic;
	PP2747 : and2 port map (X(43), Y(51), N0_51_94);
	-- signal N0_51_95 : std_logic;
	PP2748 : and2 port map (X(44), Y(51), N0_51_95);
	-- signal N0_51_96 : std_logic;
	PP2749 : and2 port map (X(45), Y(51), N0_51_96);
	-- signal N0_51_97 : std_logic;
	PP2750 : and2 port map (X(46), Y(51), N0_51_97);
	-- signal N0_51_98 : std_logic;
	PP2751 : and2 port map (X(47), Y(51), N0_51_98);
	-- signal N0_51_99 : std_logic;
	PP2752 : and2 port map (X(48), Y(51), N0_51_99);
	-- signal N0_51_100 : std_logic;
	PP2753 : and2 port map (X(49), Y(51), N0_51_100);
	-- signal N0_51_101 : std_logic;
	PP2754 : and2 port map (X(50), Y(51), N0_51_101);
	-- signal N0_51_102 : std_logic;
	PP2755 : and2 port map (X(51), Y(51), N0_51_102);
	-- signal N0_51_103 : std_logic;
	PP2756 : and2 port map ('1', Y(51), N0_51_103);
	-- signal N0_52_52 : std_logic;
	PP2757 : and2 port map (X(0), '1', N0_52_52);
	-- signal N0_52_53 : std_logic;
	PP2758 : and2 port map (X(1), '1', N0_52_53);
	-- signal N0_52_54 : std_logic;
	PP2759 : and2 port map (X(2), '1', N0_52_54);
	-- signal N0_52_55 : std_logic;
	PP2760 : and2 port map (X(3), '1', N0_52_55);
	-- signal N0_52_56 : std_logic;
	PP2761 : and2 port map (X(4), '1', N0_52_56);
	-- signal N0_52_57 : std_logic;
	PP2762 : and2 port map (X(5), '1', N0_52_57);
	-- signal N0_52_58 : std_logic;
	PP2763 : and2 port map (X(6), '1', N0_52_58);
	-- signal N0_52_59 : std_logic;
	PP2764 : and2 port map (X(7), '1', N0_52_59);
	-- signal N0_52_60 : std_logic;
	PP2765 : and2 port map (X(8), '1', N0_52_60);
	-- signal N0_52_61 : std_logic;
	PP2766 : and2 port map (X(9), '1', N0_52_61);
	-- signal N0_52_62 : std_logic;
	PP2767 : and2 port map (X(10), '1', N0_52_62);
	-- signal N0_52_63 : std_logic;
	PP2768 : and2 port map (X(11), '1', N0_52_63);
	-- signal N0_52_64 : std_logic;
	PP2769 : and2 port map (X(12), '1', N0_52_64);
	-- signal N0_52_65 : std_logic;
	PP2770 : and2 port map (X(13), '1', N0_52_65);
	-- signal N0_52_66 : std_logic;
	PP2771 : and2 port map (X(14), '1', N0_52_66);
	-- signal N0_52_67 : std_logic;
	PP2772 : and2 port map (X(15), '1', N0_52_67);
	-- signal N0_52_68 : std_logic;
	PP2773 : and2 port map (X(16), '1', N0_52_68);
	-- signal N0_52_69 : std_logic;
	PP2774 : and2 port map (X(17), '1', N0_52_69);
	-- signal N0_52_70 : std_logic;
	PP2775 : and2 port map (X(18), '1', N0_52_70);
	-- signal N0_52_71 : std_logic;
	PP2776 : and2 port map (X(19), '1', N0_52_71);
	-- signal N0_52_72 : std_logic;
	PP2777 : and2 port map (X(20), '1', N0_52_72);
	-- signal N0_52_73 : std_logic;
	PP2778 : and2 port map (X(21), '1', N0_52_73);
	-- signal N0_52_74 : std_logic;
	PP2779 : and2 port map (X(22), '1', N0_52_74);
	-- signal N0_52_75 : std_logic;
	PP2780 : and2 port map (X(23), '1', N0_52_75);
	-- signal N0_52_76 : std_logic;
	PP2781 : and2 port map (X(24), '1', N0_52_76);
	-- signal N0_52_77 : std_logic;
	PP2782 : and2 port map (X(25), '1', N0_52_77);
	-- signal N0_52_78 : std_logic;
	PP2783 : and2 port map (X(26), '1', N0_52_78);
	-- signal N0_52_79 : std_logic;
	PP2784 : and2 port map (X(27), '1', N0_52_79);
	-- signal N0_52_80 : std_logic;
	PP2785 : and2 port map (X(28), '1', N0_52_80);
	-- signal N0_52_81 : std_logic;
	PP2786 : and2 port map (X(29), '1', N0_52_81);
	-- signal N0_52_82 : std_logic;
	PP2787 : and2 port map (X(30), '1', N0_52_82);
	-- signal N0_52_83 : std_logic;
	PP2788 : and2 port map (X(31), '1', N0_52_83);
	-- signal N0_52_84 : std_logic;
	PP2789 : and2 port map (X(32), '1', N0_52_84);
	-- signal N0_52_85 : std_logic;
	PP2790 : and2 port map (X(33), '1', N0_52_85);
	-- signal N0_52_86 : std_logic;
	PP2791 : and2 port map (X(34), '1', N0_52_86);
	-- signal N0_52_87 : std_logic;
	PP2792 : and2 port map (X(35), '1', N0_52_87);
	-- signal N0_52_88 : std_logic;
	PP2793 : and2 port map (X(36), '1', N0_52_88);
	-- signal N0_52_89 : std_logic;
	PP2794 : and2 port map (X(37), '1', N0_52_89);
	-- signal N0_52_90 : std_logic;
	PP2795 : and2 port map (X(38), '1', N0_52_90);
	-- signal N0_52_91 : std_logic;
	PP2796 : and2 port map (X(39), '1', N0_52_91);
	-- signal N0_52_92 : std_logic;
	PP2797 : and2 port map (X(40), '1', N0_52_92);
	-- signal N0_52_93 : std_logic;
	PP2798 : and2 port map (X(41), '1', N0_52_93);
	-- signal N0_52_94 : std_logic;
	PP2799 : and2 port map (X(42), '1', N0_52_94);
	-- signal N0_52_95 : std_logic;
	PP2800 : and2 port map (X(43), '1', N0_52_95);
	-- signal N0_52_96 : std_logic;
	PP2801 : and2 port map (X(44), '1', N0_52_96);
	-- signal N0_52_97 : std_logic;
	PP2802 : and2 port map (X(45), '1', N0_52_97);
	-- signal N0_52_98 : std_logic;
	PP2803 : and2 port map (X(46), '1', N0_52_98);
	-- signal N0_52_99 : std_logic;
	PP2804 : and2 port map (X(47), '1', N0_52_99);
	-- signal N0_52_100 : std_logic;
	PP2805 : and2 port map (X(48), '1', N0_52_100);
	-- signal N0_52_101 : std_logic;
	PP2806 : and2 port map (X(49), '1', N0_52_101);
	-- signal N0_52_102 : std_logic;
	PP2807 : and2 port map (X(50), '1', N0_52_102);
	-- signal N0_52_103 : std_logic;
	PP2808 : and2 port map (X(51), '1', N0_52_103);
	-- signal N0_52_104 : std_logic;
	PP2809 : and2 port map ('1', '1', N0_52_104);

-- PP Reduction
	-- Elements from matrix 0 
	-- Elements from matrix 1 
-- In matrix 1 adding HA to column 36 
	-- signal N2_0_36 : std_logic;
	-- signal N2_1_37 : std_logic;
	HA1 : half_adder port map (N0_0_36,N0_1_36,N2_0_36,N2_1_37);
-- In matrix 1 adding FA to column 37 
	-- signal N2_0_37 : std_logic;
	-- signal N2_1_38 : std_logic;
	FA1 : full_adder port map (N0_0_37,N0_1_37,N0_2_37,N2_0_37,N2_1_38);
-- In matrix 1 adding HA to column 37 
	-- signal N2_2_37 : std_logic;
	-- signal N2_3_38 : std_logic;
	HA2 : half_adder port map (N0_3_37,N0_4_37,N2_2_37,N2_3_38);
-- In matrix 1 adding FA to column 38 
	-- signal N2_0_38 : std_logic;
	-- signal N2_1_39 : std_logic;
	FA2 : full_adder port map (N0_0_38,N0_1_38,N0_2_38,N2_0_38,N2_1_39);
-- In matrix 1 adding FA to column 38 
	-- signal N2_2_38 : std_logic;
	-- signal N2_3_39 : std_logic;
	FA3 : full_adder port map (N0_3_38,N0_4_38,N0_5_38,N2_2_38,N2_3_39);
-- In matrix 1 adding HA to column 38 
	-- signal N2_4_38 : std_logic;
	-- signal N2_5_39 : std_logic;
	HA3 : half_adder port map (N0_6_38,N0_7_38,N2_4_38,N2_5_39);
-- In matrix 1 adding FA to column 39 
	-- signal N2_0_39 : std_logic;
	-- signal N2_1_40 : std_logic;
	FA4 : full_adder port map (N0_0_39,N0_1_39,N0_2_39,N2_0_39,N2_1_40);
-- In matrix 1 adding FA to column 39 
	-- signal N2_2_39 : std_logic;
	-- signal N2_3_40 : std_logic;
	FA5 : full_adder port map (N0_3_39,N0_4_39,N0_5_39,N2_2_39,N2_3_40);
-- In matrix 1 adding FA to column 39 
	-- signal N2_4_39 : std_logic;
	-- signal N2_5_40 : std_logic;
	FA6 : full_adder port map (N0_6_39,N0_7_39,N0_8_39,N2_4_39,N2_5_40);
-- In matrix 1 adding HA to column 39 
	-- signal N2_6_39 : std_logic;
	-- signal N2_7_40 : std_logic;
	HA4 : half_adder port map (N0_9_39,N0_10_39,N2_6_39,N2_7_40);
-- In matrix 1 adding FA to column 40 
	-- signal N2_0_40 : std_logic;
	-- signal N2_1_41 : std_logic;
	FA7 : full_adder port map (N0_0_40,N0_1_40,N0_2_40,N2_0_40,N2_1_41);
-- In matrix 1 adding FA to column 40 
	-- signal N2_2_40 : std_logic;
	-- signal N2_3_41 : std_logic;
	FA8 : full_adder port map (N0_3_40,N0_4_40,N0_5_40,N2_2_40,N2_3_41);
-- In matrix 1 adding FA to column 40 
	-- signal N2_4_40 : std_logic;
	-- signal N2_5_41 : std_logic;
	FA9 : full_adder port map (N0_6_40,N0_7_40,N0_8_40,N2_4_40,N2_5_41);
-- In matrix 1 adding FA to column 40 
	-- signal N2_6_40 : std_logic;
	-- signal N2_7_41 : std_logic;
	FA10 : full_adder port map (N0_9_40,N0_10_40,N0_11_40,N2_6_40,N2_7_41);
-- In matrix 1 adding HA to column 40 
	-- signal N2_8_40 : std_logic;
	-- signal N2_9_41 : std_logic;
	HA5 : half_adder port map (N0_12_40,N0_13_40,N2_8_40,N2_9_41);
-- In matrix 1 adding FA to column 41 
	-- signal N2_0_41 : std_logic;
	-- signal N2_1_42 : std_logic;
	FA11 : full_adder port map (N0_0_41,N0_1_41,N0_2_41,N2_0_41,N2_1_42);
-- In matrix 1 adding FA to column 41 
	-- signal N2_2_41 : std_logic;
	-- signal N2_3_42 : std_logic;
	FA12 : full_adder port map (N0_3_41,N0_4_41,N0_5_41,N2_2_41,N2_3_42);
-- In matrix 1 adding FA to column 41 
	-- signal N2_4_41 : std_logic;
	-- signal N2_5_42 : std_logic;
	FA13 : full_adder port map (N0_6_41,N0_7_41,N0_8_41,N2_4_41,N2_5_42);
-- In matrix 1 adding FA to column 41 
	-- signal N2_6_41 : std_logic;
	-- signal N2_7_42 : std_logic;
	FA14 : full_adder port map (N0_9_41,N0_10_41,N0_11_41,N2_6_41,N2_7_42);
-- In matrix 1 adding FA to column 41 
	-- signal N2_8_41 : std_logic;
	-- signal N2_9_42 : std_logic;
	FA15 : full_adder port map (N0_12_41,N0_13_41,N0_14_41,N2_8_41,N2_9_42);
-- In matrix 1 adding HA to column 41 
	-- signal N2_10_41 : std_logic;
	-- signal N2_11_42 : std_logic;
	HA6 : half_adder port map (N0_15_41,N0_16_41,N2_10_41,N2_11_42);
-- In matrix 1 adding FA to column 42 
	-- signal N2_0_42 : std_logic;
	-- signal N2_1_43 : std_logic;
	FA16 : full_adder port map (N0_0_42,N0_1_42,N0_2_42,N2_0_42,N2_1_43);
-- In matrix 1 adding FA to column 42 
	-- signal N2_2_42 : std_logic;
	-- signal N2_3_43 : std_logic;
	FA17 : full_adder port map (N0_3_42,N0_4_42,N0_5_42,N2_2_42,N2_3_43);
-- In matrix 1 adding FA to column 42 
	-- signal N2_4_42 : std_logic;
	-- signal N2_5_43 : std_logic;
	FA18 : full_adder port map (N0_6_42,N0_7_42,N0_8_42,N2_4_42,N2_5_43);
-- In matrix 1 adding FA to column 42 
	-- signal N2_6_42 : std_logic;
	-- signal N2_7_43 : std_logic;
	FA19 : full_adder port map (N0_9_42,N0_10_42,N0_11_42,N2_6_42,N2_7_43);
-- In matrix 1 adding FA to column 42 
	-- signal N2_8_42 : std_logic;
	-- signal N2_9_43 : std_logic;
	FA20 : full_adder port map (N0_12_42,N0_13_42,N0_14_42,N2_8_42,N2_9_43);
-- In matrix 1 adding FA to column 42 
	-- signal N2_10_42 : std_logic;
	-- signal N2_11_43 : std_logic;
	FA21 : full_adder port map (N0_15_42,N0_16_42,N0_17_42,N2_10_42,N2_11_43);
-- In matrix 1 adding HA to column 42 
	-- signal N2_12_42 : std_logic;
	-- signal N2_13_43 : std_logic;
	HA7 : half_adder port map (N0_18_42,N0_19_42,N2_12_42,N2_13_43);
-- In matrix 1 adding FA to column 43 
	-- signal N2_0_43 : std_logic;
	-- signal N2_1_44 : std_logic;
	FA22 : full_adder port map (N0_0_43,N0_1_43,N0_2_43,N2_0_43,N2_1_44);
-- In matrix 1 adding FA to column 43 
	-- signal N2_2_43 : std_logic;
	-- signal N2_3_44 : std_logic;
	FA23 : full_adder port map (N0_3_43,N0_4_43,N0_5_43,N2_2_43,N2_3_44);
-- In matrix 1 adding FA to column 43 
	-- signal N2_4_43 : std_logic;
	-- signal N2_5_44 : std_logic;
	FA24 : full_adder port map (N0_6_43,N0_7_43,N0_8_43,N2_4_43,N2_5_44);
-- In matrix 1 adding FA to column 43 
	-- signal N2_6_43 : std_logic;
	-- signal N2_7_44 : std_logic;
	FA25 : full_adder port map (N0_9_43,N0_10_43,N0_11_43,N2_6_43,N2_7_44);
-- In matrix 1 adding FA to column 43 
	-- signal N2_8_43 : std_logic;
	-- signal N2_9_44 : std_logic;
	FA26 : full_adder port map (N0_12_43,N0_13_43,N0_14_43,N2_8_43,N2_9_44);
-- In matrix 1 adding FA to column 43 
	-- signal N2_10_43 : std_logic;
	-- signal N2_11_44 : std_logic;
	FA27 : full_adder port map (N0_15_43,N0_16_43,N0_17_43,N2_10_43,N2_11_44);
-- In matrix 1 adding FA to column 43 
	-- signal N2_12_43 : std_logic;
	-- signal N2_13_44 : std_logic;
	FA28 : full_adder port map (N0_18_43,N0_19_43,N0_20_43,N2_12_43,N2_13_44);
-- In matrix 1 adding HA to column 43 
	-- signal N2_14_43 : std_logic;
	-- signal N2_15_44 : std_logic;
	HA8 : half_adder port map (N0_21_43,N0_22_43,N2_14_43,N2_15_44);
-- In matrix 1 adding FA to column 44 
	-- signal N2_0_44 : std_logic;
	-- signal N2_1_45 : std_logic;
	FA29 : full_adder port map (N0_0_44,N0_1_44,N0_2_44,N2_0_44,N2_1_45);
-- In matrix 1 adding FA to column 44 
	-- signal N2_2_44 : std_logic;
	-- signal N2_3_45 : std_logic;
	FA30 : full_adder port map (N0_3_44,N0_4_44,N0_5_44,N2_2_44,N2_3_45);
-- In matrix 1 adding FA to column 44 
	-- signal N2_4_44 : std_logic;
	-- signal N2_5_45 : std_logic;
	FA31 : full_adder port map (N0_6_44,N0_7_44,N0_8_44,N2_4_44,N2_5_45);
-- In matrix 1 adding FA to column 44 
	-- signal N2_6_44 : std_logic;
	-- signal N2_7_45 : std_logic;
	FA32 : full_adder port map (N0_9_44,N0_10_44,N0_11_44,N2_6_44,N2_7_45);
-- In matrix 1 adding FA to column 44 
	-- signal N2_8_44 : std_logic;
	-- signal N2_9_45 : std_logic;
	FA33 : full_adder port map (N0_12_44,N0_13_44,N0_14_44,N2_8_44,N2_9_45);
-- In matrix 1 adding FA to column 44 
	-- signal N2_10_44 : std_logic;
	-- signal N2_11_45 : std_logic;
	FA34 : full_adder port map (N0_15_44,N0_16_44,N0_17_44,N2_10_44,N2_11_45);
-- In matrix 1 adding FA to column 44 
	-- signal N2_12_44 : std_logic;
	-- signal N2_13_45 : std_logic;
	FA35 : full_adder port map (N0_18_44,N0_19_44,N0_20_44,N2_12_44,N2_13_45);
-- In matrix 1 adding FA to column 44 
	-- signal N2_14_44 : std_logic;
	-- signal N2_15_45 : std_logic;
	FA36 : full_adder port map (N0_21_44,N0_22_44,N0_23_44,N2_14_44,N2_15_45);
-- In matrix 1 adding HA to column 44 
	-- signal N2_16_44 : std_logic;
	-- signal N2_17_45 : std_logic;
	HA9 : half_adder port map (N0_24_44,N0_25_44,N2_16_44,N2_17_45);
-- In matrix 1 adding FA to column 45 
	-- signal N2_0_45 : std_logic;
	-- signal N2_1_46 : std_logic;
	FA37 : full_adder port map (N0_0_45,N0_1_45,N0_2_45,N2_0_45,N2_1_46);
-- In matrix 1 adding FA to column 45 
	-- signal N2_2_45 : std_logic;
	-- signal N2_3_46 : std_logic;
	FA38 : full_adder port map (N0_3_45,N0_4_45,N0_5_45,N2_2_45,N2_3_46);
-- In matrix 1 adding FA to column 45 
	-- signal N2_4_45 : std_logic;
	-- signal N2_5_46 : std_logic;
	FA39 : full_adder port map (N0_6_45,N0_7_45,N0_8_45,N2_4_45,N2_5_46);
-- In matrix 1 adding FA to column 45 
	-- signal N2_6_45 : std_logic;
	-- signal N2_7_46 : std_logic;
	FA40 : full_adder port map (N0_9_45,N0_10_45,N0_11_45,N2_6_45,N2_7_46);
-- In matrix 1 adding FA to column 45 
	-- signal N2_8_45 : std_logic;
	-- signal N2_9_46 : std_logic;
	FA41 : full_adder port map (N0_12_45,N0_13_45,N0_14_45,N2_8_45,N2_9_46);
-- In matrix 1 adding FA to column 45 
	-- signal N2_10_45 : std_logic;
	-- signal N2_11_46 : std_logic;
	FA42 : full_adder port map (N0_15_45,N0_16_45,N0_17_45,N2_10_45,N2_11_46);
-- In matrix 1 adding FA to column 45 
	-- signal N2_12_45 : std_logic;
	-- signal N2_13_46 : std_logic;
	FA43 : full_adder port map (N0_18_45,N0_19_45,N0_20_45,N2_12_45,N2_13_46);
-- In matrix 1 adding FA to column 45 
	-- signal N2_14_45 : std_logic;
	-- signal N2_15_46 : std_logic;
	FA44 : full_adder port map (N0_21_45,N0_22_45,N0_23_45,N2_14_45,N2_15_46);
-- In matrix 1 adding FA to column 45 
	-- signal N2_16_45 : std_logic;
	-- signal N2_17_46 : std_logic;
	FA45 : full_adder port map (N0_24_45,N0_25_45,N0_26_45,N2_16_45,N2_17_46);
-- In matrix 1 adding HA to column 45 
	-- signal N2_18_45 : std_logic;
	-- signal N2_19_46 : std_logic;
	HA10 : half_adder port map (N0_27_45,N0_28_45,N2_18_45,N2_19_46);
-- In matrix 1 adding FA to column 46 
	-- signal N2_0_46 : std_logic;
	-- signal N2_1_47 : std_logic;
	FA46 : full_adder port map (N0_0_46,N0_1_46,N0_2_46,N2_0_46,N2_1_47);
-- In matrix 1 adding FA to column 46 
	-- signal N2_2_46 : std_logic;
	-- signal N2_3_47 : std_logic;
	FA47 : full_adder port map (N0_3_46,N0_4_46,N0_5_46,N2_2_46,N2_3_47);
-- In matrix 1 adding FA to column 46 
	-- signal N2_4_46 : std_logic;
	-- signal N2_5_47 : std_logic;
	FA48 : full_adder port map (N0_6_46,N0_7_46,N0_8_46,N2_4_46,N2_5_47);
-- In matrix 1 adding FA to column 46 
	-- signal N2_6_46 : std_logic;
	-- signal N2_7_47 : std_logic;
	FA49 : full_adder port map (N0_9_46,N0_10_46,N0_11_46,N2_6_46,N2_7_47);
-- In matrix 1 adding FA to column 46 
	-- signal N2_8_46 : std_logic;
	-- signal N2_9_47 : std_logic;
	FA50 : full_adder port map (N0_12_46,N0_13_46,N0_14_46,N2_8_46,N2_9_47);
-- In matrix 1 adding FA to column 46 
	-- signal N2_10_46 : std_logic;
	-- signal N2_11_47 : std_logic;
	FA51 : full_adder port map (N0_15_46,N0_16_46,N0_17_46,N2_10_46,N2_11_47);
-- In matrix 1 adding FA to column 46 
	-- signal N2_12_46 : std_logic;
	-- signal N2_13_47 : std_logic;
	FA52 : full_adder port map (N0_18_46,N0_19_46,N0_20_46,N2_12_46,N2_13_47);
-- In matrix 1 adding FA to column 46 
	-- signal N2_14_46 : std_logic;
	-- signal N2_15_47 : std_logic;
	FA53 : full_adder port map (N0_21_46,N0_22_46,N0_23_46,N2_14_46,N2_15_47);
-- In matrix 1 adding FA to column 46 
	-- signal N2_16_46 : std_logic;
	-- signal N2_17_47 : std_logic;
	FA54 : full_adder port map (N0_24_46,N0_25_46,N0_26_46,N2_16_46,N2_17_47);
-- In matrix 1 adding FA to column 46 
	-- signal N2_18_46 : std_logic;
	-- signal N2_19_47 : std_logic;
	FA55 : full_adder port map (N0_27_46,N0_28_46,N0_29_46,N2_18_46,N2_19_47);
-- In matrix 1 adding HA to column 46 
	-- signal N2_20_46 : std_logic;
	-- signal N2_21_47 : std_logic;
	HA11 : half_adder port map (N0_30_46,N0_31_46,N2_20_46,N2_21_47);
-- In matrix 1 adding FA to column 47 
	-- signal N2_0_47 : std_logic;
	-- signal N2_1_48 : std_logic;
	FA56 : full_adder port map (N0_0_47,N0_1_47,N0_2_47,N2_0_47,N2_1_48);
-- In matrix 1 adding FA to column 47 
	-- signal N2_2_47 : std_logic;
	-- signal N2_3_48 : std_logic;
	FA57 : full_adder port map (N0_3_47,N0_4_47,N0_5_47,N2_2_47,N2_3_48);
-- In matrix 1 adding FA to column 47 
	-- signal N2_4_47 : std_logic;
	-- signal N2_5_48 : std_logic;
	FA58 : full_adder port map (N0_6_47,N0_7_47,N0_8_47,N2_4_47,N2_5_48);
-- In matrix 1 adding FA to column 47 
	-- signal N2_6_47 : std_logic;
	-- signal N2_7_48 : std_logic;
	FA59 : full_adder port map (N0_9_47,N0_10_47,N0_11_47,N2_6_47,N2_7_48);
-- In matrix 1 adding FA to column 47 
	-- signal N2_8_47 : std_logic;
	-- signal N2_9_48 : std_logic;
	FA60 : full_adder port map (N0_12_47,N0_13_47,N0_14_47,N2_8_47,N2_9_48);
-- In matrix 1 adding FA to column 47 
	-- signal N2_10_47 : std_logic;
	-- signal N2_11_48 : std_logic;
	FA61 : full_adder port map (N0_15_47,N0_16_47,N0_17_47,N2_10_47,N2_11_48);
-- In matrix 1 adding FA to column 47 
	-- signal N2_12_47 : std_logic;
	-- signal N2_13_48 : std_logic;
	FA62 : full_adder port map (N0_18_47,N0_19_47,N0_20_47,N2_12_47,N2_13_48);
-- In matrix 1 adding FA to column 47 
	-- signal N2_14_47 : std_logic;
	-- signal N2_15_48 : std_logic;
	FA63 : full_adder port map (N0_21_47,N0_22_47,N0_23_47,N2_14_47,N2_15_48);
-- In matrix 1 adding FA to column 47 
	-- signal N2_16_47 : std_logic;
	-- signal N2_17_48 : std_logic;
	FA64 : full_adder port map (N0_24_47,N0_25_47,N0_26_47,N2_16_47,N2_17_48);
-- In matrix 1 adding FA to column 47 
	-- signal N2_18_47 : std_logic;
	-- signal N2_19_48 : std_logic;
	FA65 : full_adder port map (N0_27_47,N0_28_47,N0_29_47,N2_18_47,N2_19_48);
-- In matrix 1 adding FA to column 47 
	-- signal N2_20_47 : std_logic;
	-- signal N2_21_48 : std_logic;
	FA66 : full_adder port map (N0_30_47,N0_31_47,N0_32_47,N2_20_47,N2_21_48);
-- In matrix 1 adding HA to column 47 
	-- signal N2_22_47 : std_logic;
	-- signal N2_23_48 : std_logic;
	HA12 : half_adder port map (N0_33_47,N0_34_47,N2_22_47,N2_23_48);
-- In matrix 1 adding FA to column 48 
	-- signal N2_0_48 : std_logic;
	-- signal N2_1_49 : std_logic;
	FA67 : full_adder port map (N0_0_48,N0_1_48,N0_2_48,N2_0_48,N2_1_49);
-- In matrix 1 adding FA to column 48 
	-- signal N2_2_48 : std_logic;
	-- signal N2_3_49 : std_logic;
	FA68 : full_adder port map (N0_3_48,N0_4_48,N0_5_48,N2_2_48,N2_3_49);
-- In matrix 1 adding FA to column 48 
	-- signal N2_4_48 : std_logic;
	-- signal N2_5_49 : std_logic;
	FA69 : full_adder port map (N0_6_48,N0_7_48,N0_8_48,N2_4_48,N2_5_49);
-- In matrix 1 adding FA to column 48 
	-- signal N2_6_48 : std_logic;
	-- signal N2_7_49 : std_logic;
	FA70 : full_adder port map (N0_9_48,N0_10_48,N0_11_48,N2_6_48,N2_7_49);
-- In matrix 1 adding FA to column 48 
	-- signal N2_8_48 : std_logic;
	-- signal N2_9_49 : std_logic;
	FA71 : full_adder port map (N0_12_48,N0_13_48,N0_14_48,N2_8_48,N2_9_49);
-- In matrix 1 adding FA to column 48 
	-- signal N2_10_48 : std_logic;
	-- signal N2_11_49 : std_logic;
	FA72 : full_adder port map (N0_15_48,N0_16_48,N0_17_48,N2_10_48,N2_11_49);
-- In matrix 1 adding FA to column 48 
	-- signal N2_12_48 : std_logic;
	-- signal N2_13_49 : std_logic;
	FA73 : full_adder port map (N0_18_48,N0_19_48,N0_20_48,N2_12_48,N2_13_49);
-- In matrix 1 adding FA to column 48 
	-- signal N2_14_48 : std_logic;
	-- signal N2_15_49 : std_logic;
	FA74 : full_adder port map (N0_21_48,N0_22_48,N0_23_48,N2_14_48,N2_15_49);
-- In matrix 1 adding FA to column 48 
	-- signal N2_16_48 : std_logic;
	-- signal N2_17_49 : std_logic;
	FA75 : full_adder port map (N0_24_48,N0_25_48,N0_26_48,N2_16_48,N2_17_49);
-- In matrix 1 adding FA to column 48 
	-- signal N2_18_48 : std_logic;
	-- signal N2_19_49 : std_logic;
	FA76 : full_adder port map (N0_27_48,N0_28_48,N0_29_48,N2_18_48,N2_19_49);
-- In matrix 1 adding FA to column 48 
	-- signal N2_20_48 : std_logic;
	-- signal N2_21_49 : std_logic;
	FA77 : full_adder port map (N0_30_48,N0_31_48,N0_32_48,N2_20_48,N2_21_49);
-- In matrix 1 adding FA to column 48 
	-- signal N2_22_48 : std_logic;
	-- signal N2_23_49 : std_logic;
	FA78 : full_adder port map (N0_33_48,N0_34_48,N0_35_48,N2_22_48,N2_23_49);
-- In matrix 1 adding HA to column 48 
	-- signal N2_24_48 : std_logic;
	-- signal N2_25_49 : std_logic;
	HA13 : half_adder port map (N0_36_48,N0_37_48,N2_24_48,N2_25_49);
-- In matrix 1 adding FA to column 49 
	-- signal N2_0_49 : std_logic;
	-- signal N2_1_50 : std_logic;
	FA79 : full_adder port map (N0_0_49,N0_1_49,N0_2_49,N2_0_49,N2_1_50);
-- In matrix 1 adding FA to column 49 
	-- signal N2_2_49 : std_logic;
	-- signal N2_3_50 : std_logic;
	FA80 : full_adder port map (N0_3_49,N0_4_49,N0_5_49,N2_2_49,N2_3_50);
-- In matrix 1 adding FA to column 49 
	-- signal N2_4_49 : std_logic;
	-- signal N2_5_50 : std_logic;
	FA81 : full_adder port map (N0_6_49,N0_7_49,N0_8_49,N2_4_49,N2_5_50);
-- In matrix 1 adding FA to column 49 
	-- signal N2_6_49 : std_logic;
	-- signal N2_7_50 : std_logic;
	FA82 : full_adder port map (N0_9_49,N0_10_49,N0_11_49,N2_6_49,N2_7_50);
-- In matrix 1 adding FA to column 49 
	-- signal N2_8_49 : std_logic;
	-- signal N2_9_50 : std_logic;
	FA83 : full_adder port map (N0_12_49,N0_13_49,N0_14_49,N2_8_49,N2_9_50);
-- In matrix 1 adding FA to column 49 
	-- signal N2_10_49 : std_logic;
	-- signal N2_11_50 : std_logic;
	FA84 : full_adder port map (N0_15_49,N0_16_49,N0_17_49,N2_10_49,N2_11_50);
-- In matrix 1 adding FA to column 49 
	-- signal N2_12_49 : std_logic;
	-- signal N2_13_50 : std_logic;
	FA85 : full_adder port map (N0_18_49,N0_19_49,N0_20_49,N2_12_49,N2_13_50);
-- In matrix 1 adding FA to column 49 
	-- signal N2_14_49 : std_logic;
	-- signal N2_15_50 : std_logic;
	FA86 : full_adder port map (N0_21_49,N0_22_49,N0_23_49,N2_14_49,N2_15_50);
-- In matrix 1 adding FA to column 49 
	-- signal N2_16_49 : std_logic;
	-- signal N2_17_50 : std_logic;
	FA87 : full_adder port map (N0_24_49,N0_25_49,N0_26_49,N2_16_49,N2_17_50);
-- In matrix 1 adding FA to column 49 
	-- signal N2_18_49 : std_logic;
	-- signal N2_19_50 : std_logic;
	FA88 : full_adder port map (N0_27_49,N0_28_49,N0_29_49,N2_18_49,N2_19_50);
-- In matrix 1 adding FA to column 49 
	-- signal N2_20_49 : std_logic;
	-- signal N2_21_50 : std_logic;
	FA89 : full_adder port map (N0_30_49,N0_31_49,N0_32_49,N2_20_49,N2_21_50);
-- In matrix 1 adding FA to column 49 
	-- signal N2_22_49 : std_logic;
	-- signal N2_23_50 : std_logic;
	FA90 : full_adder port map (N0_33_49,N0_34_49,N0_35_49,N2_22_49,N2_23_50);
-- In matrix 1 adding FA to column 49 
	-- signal N2_24_49 : std_logic;
	-- signal N2_25_50 : std_logic;
	FA91 : full_adder port map (N0_36_49,N0_37_49,N0_38_49,N2_24_49,N2_25_50);
-- In matrix 1 adding HA to column 49 
	-- signal N2_26_49 : std_logic;
	-- signal N2_27_50 : std_logic;
	HA14 : half_adder port map (N0_39_49,N0_40_49,N2_26_49,N2_27_50);
-- In matrix 1 adding FA to column 50 
	-- signal N2_0_50 : std_logic;
	-- signal N2_1_51 : std_logic;
	FA92 : full_adder port map (N0_0_50,N0_1_50,N0_2_50,N2_0_50,N2_1_51);
-- In matrix 1 adding FA to column 50 
	-- signal N2_2_50 : std_logic;
	-- signal N2_3_51 : std_logic;
	FA93 : full_adder port map (N0_3_50,N0_4_50,N0_5_50,N2_2_50,N2_3_51);
-- In matrix 1 adding FA to column 50 
	-- signal N2_4_50 : std_logic;
	-- signal N2_5_51 : std_logic;
	FA94 : full_adder port map (N0_6_50,N0_7_50,N0_8_50,N2_4_50,N2_5_51);
-- In matrix 1 adding FA to column 50 
	-- signal N2_6_50 : std_logic;
	-- signal N2_7_51 : std_logic;
	FA95 : full_adder port map (N0_9_50,N0_10_50,N0_11_50,N2_6_50,N2_7_51);
-- In matrix 1 adding FA to column 50 
	-- signal N2_8_50 : std_logic;
	-- signal N2_9_51 : std_logic;
	FA96 : full_adder port map (N0_12_50,N0_13_50,N0_14_50,N2_8_50,N2_9_51);
-- In matrix 1 adding FA to column 50 
	-- signal N2_10_50 : std_logic;
	-- signal N2_11_51 : std_logic;
	FA97 : full_adder port map (N0_15_50,N0_16_50,N0_17_50,N2_10_50,N2_11_51);
-- In matrix 1 adding FA to column 50 
	-- signal N2_12_50 : std_logic;
	-- signal N2_13_51 : std_logic;
	FA98 : full_adder port map (N0_18_50,N0_19_50,N0_20_50,N2_12_50,N2_13_51);
-- In matrix 1 adding FA to column 50 
	-- signal N2_14_50 : std_logic;
	-- signal N2_15_51 : std_logic;
	FA99 : full_adder port map (N0_21_50,N0_22_50,N0_23_50,N2_14_50,N2_15_51);
-- In matrix 1 adding FA to column 50 
	-- signal N2_16_50 : std_logic;
	-- signal N2_17_51 : std_logic;
	FA100 : full_adder port map (N0_24_50,N0_25_50,N0_26_50,N2_16_50,N2_17_51);
-- In matrix 1 adding FA to column 50 
	-- signal N2_18_50 : std_logic;
	-- signal N2_19_51 : std_logic;
	FA101 : full_adder port map (N0_27_50,N0_28_50,N0_29_50,N2_18_50,N2_19_51);
-- In matrix 1 adding FA to column 50 
	-- signal N2_20_50 : std_logic;
	-- signal N2_21_51 : std_logic;
	FA102 : full_adder port map (N0_30_50,N0_31_50,N0_32_50,N2_20_50,N2_21_51);
-- In matrix 1 adding FA to column 50 
	-- signal N2_22_50 : std_logic;
	-- signal N2_23_51 : std_logic;
	FA103 : full_adder port map (N0_33_50,N0_34_50,N0_35_50,N2_22_50,N2_23_51);
-- In matrix 1 adding FA to column 50 
	-- signal N2_24_50 : std_logic;
	-- signal N2_25_51 : std_logic;
	FA104 : full_adder port map (N0_36_50,N0_37_50,N0_38_50,N2_24_50,N2_25_51);
-- In matrix 1 adding FA to column 50 
	-- signal N2_26_50 : std_logic;
	-- signal N2_27_51 : std_logic;
	FA105 : full_adder port map (N0_39_50,N0_40_50,N0_41_50,N2_26_50,N2_27_51);
-- In matrix 1 adding HA to column 50 
	-- signal N2_28_50 : std_logic;
	-- signal N2_29_51 : std_logic;
	HA15 : half_adder port map (N0_42_50,N0_43_50,N2_28_50,N2_29_51);
-- In matrix 1 adding FA to column 51 
	-- signal N2_0_51 : std_logic;
	-- signal N2_1_52 : std_logic;
	FA106 : full_adder port map (N0_0_51,N0_1_51,N0_2_51,N2_0_51,N2_1_52);
-- In matrix 1 adding FA to column 51 
	-- signal N2_2_51 : std_logic;
	-- signal N2_3_52 : std_logic;
	FA107 : full_adder port map (N0_3_51,N0_4_51,N0_5_51,N2_2_51,N2_3_52);
-- In matrix 1 adding FA to column 51 
	-- signal N2_4_51 : std_logic;
	-- signal N2_5_52 : std_logic;
	FA108 : full_adder port map (N0_6_51,N0_7_51,N0_8_51,N2_4_51,N2_5_52);
-- In matrix 1 adding FA to column 51 
	-- signal N2_6_51 : std_logic;
	-- signal N2_7_52 : std_logic;
	FA109 : full_adder port map (N0_9_51,N0_10_51,N0_11_51,N2_6_51,N2_7_52);
-- In matrix 1 adding FA to column 51 
	-- signal N2_8_51 : std_logic;
	-- signal N2_9_52 : std_logic;
	FA110 : full_adder port map (N0_12_51,N0_13_51,N0_14_51,N2_8_51,N2_9_52);
-- In matrix 1 adding FA to column 51 
	-- signal N2_10_51 : std_logic;
	-- signal N2_11_52 : std_logic;
	FA111 : full_adder port map (N0_15_51,N0_16_51,N0_17_51,N2_10_51,N2_11_52);
-- In matrix 1 adding FA to column 51 
	-- signal N2_12_51 : std_logic;
	-- signal N2_13_52 : std_logic;
	FA112 : full_adder port map (N0_18_51,N0_19_51,N0_20_51,N2_12_51,N2_13_52);
-- In matrix 1 adding FA to column 51 
	-- signal N2_14_51 : std_logic;
	-- signal N2_15_52 : std_logic;
	FA113 : full_adder port map (N0_21_51,N0_22_51,N0_23_51,N2_14_51,N2_15_52);
-- In matrix 1 adding FA to column 51 
	-- signal N2_16_51 : std_logic;
	-- signal N2_17_52 : std_logic;
	FA114 : full_adder port map (N0_24_51,N0_25_51,N0_26_51,N2_16_51,N2_17_52);
-- In matrix 1 adding FA to column 51 
	-- signal N2_18_51 : std_logic;
	-- signal N2_19_52 : std_logic;
	FA115 : full_adder port map (N0_27_51,N0_28_51,N0_29_51,N2_18_51,N2_19_52);
-- In matrix 1 adding FA to column 51 
	-- signal N2_20_51 : std_logic;
	-- signal N2_21_52 : std_logic;
	FA116 : full_adder port map (N0_30_51,N0_31_51,N0_32_51,N2_20_51,N2_21_52);
-- In matrix 1 adding FA to column 51 
	-- signal N2_22_51 : std_logic;
	-- signal N2_23_52 : std_logic;
	FA117 : full_adder port map (N0_33_51,N0_34_51,N0_35_51,N2_22_51,N2_23_52);
-- In matrix 1 adding FA to column 51 
	-- signal N2_24_51 : std_logic;
	-- signal N2_25_52 : std_logic;
	FA118 : full_adder port map (N0_36_51,N0_37_51,N0_38_51,N2_24_51,N2_25_52);
-- In matrix 1 adding FA to column 51 
	-- signal N2_26_51 : std_logic;
	-- signal N2_27_52 : std_logic;
	FA119 : full_adder port map (N0_39_51,N0_40_51,N0_41_51,N2_26_51,N2_27_52);
-- In matrix 1 adding FA to column 51 
	-- signal N2_28_51 : std_logic;
	-- signal N2_29_52 : std_logic;
	FA120 : full_adder port map (N0_42_51,N0_43_51,N0_44_51,N2_28_51,N2_29_52);
-- In matrix 1 adding HA to column 51 
	-- signal N2_30_51 : std_logic;
	-- signal N2_31_52 : std_logic;
	HA16 : half_adder port map (N0_45_51,N0_46_51,N2_30_51,N2_31_52);
-- In matrix 1 adding FA to column 52 
	-- signal N2_0_52 : std_logic;
	-- signal N2_1_53 : std_logic;
	FA121 : full_adder port map (N0_0_52,N0_1_52,N0_2_52,N2_0_52,N2_1_53);
-- In matrix 1 adding FA to column 52 
	-- signal N2_2_52 : std_logic;
	-- signal N2_3_53 : std_logic;
	FA122 : full_adder port map (N0_3_52,N0_4_52,N0_5_52,N2_2_52,N2_3_53);
-- In matrix 1 adding FA to column 52 
	-- signal N2_4_52 : std_logic;
	-- signal N2_5_53 : std_logic;
	FA123 : full_adder port map (N0_6_52,N0_7_52,N0_8_52,N2_4_52,N2_5_53);
-- In matrix 1 adding FA to column 52 
	-- signal N2_6_52 : std_logic;
	-- signal N2_7_53 : std_logic;
	FA124 : full_adder port map (N0_9_52,N0_10_52,N0_11_52,N2_6_52,N2_7_53);
-- In matrix 1 adding FA to column 52 
	-- signal N2_8_52 : std_logic;
	-- signal N2_9_53 : std_logic;
	FA125 : full_adder port map (N0_12_52,N0_13_52,N0_14_52,N2_8_52,N2_9_53);
-- In matrix 1 adding FA to column 52 
	-- signal N2_10_52 : std_logic;
	-- signal N2_11_53 : std_logic;
	FA126 : full_adder port map (N0_15_52,N0_16_52,N0_17_52,N2_10_52,N2_11_53);
-- In matrix 1 adding FA to column 52 
	-- signal N2_12_52 : std_logic;
	-- signal N2_13_53 : std_logic;
	FA127 : full_adder port map (N0_18_52,N0_19_52,N0_20_52,N2_12_52,N2_13_53);
-- In matrix 1 adding FA to column 52 
	-- signal N2_14_52 : std_logic;
	-- signal N2_15_53 : std_logic;
	FA128 : full_adder port map (N0_21_52,N0_22_52,N0_23_52,N2_14_52,N2_15_53);
-- In matrix 1 adding FA to column 52 
	-- signal N2_16_52 : std_logic;
	-- signal N2_17_53 : std_logic;
	FA129 : full_adder port map (N0_24_52,N0_25_52,N0_26_52,N2_16_52,N2_17_53);
-- In matrix 1 adding FA to column 52 
	-- signal N2_18_52 : std_logic;
	-- signal N2_19_53 : std_logic;
	FA130 : full_adder port map (N0_27_52,N0_28_52,N0_29_52,N2_18_52,N2_19_53);
-- In matrix 1 adding FA to column 52 
	-- signal N2_20_52 : std_logic;
	-- signal N2_21_53 : std_logic;
	FA131 : full_adder port map (N0_30_52,N0_31_52,N0_32_52,N2_20_52,N2_21_53);
-- In matrix 1 adding FA to column 52 
	-- signal N2_22_52 : std_logic;
	-- signal N2_23_53 : std_logic;
	FA132 : full_adder port map (N0_33_52,N0_34_52,N0_35_52,N2_22_52,N2_23_53);
-- In matrix 1 adding FA to column 52 
	-- signal N2_24_52 : std_logic;
	-- signal N2_25_53 : std_logic;
	FA133 : full_adder port map (N0_36_52,N0_37_52,N0_38_52,N2_24_52,N2_25_53);
-- In matrix 1 adding FA to column 52 
	-- signal N2_26_52 : std_logic;
	-- signal N2_27_53 : std_logic;
	FA134 : full_adder port map (N0_39_52,N0_40_52,N0_41_52,N2_26_52,N2_27_53);
-- In matrix 1 adding FA to column 52 
	-- signal N2_28_52 : std_logic;
	-- signal N2_29_53 : std_logic;
	FA135 : full_adder port map (N0_42_52,N0_43_52,N0_44_52,N2_28_52,N2_29_53);
-- In matrix 1 adding FA to column 52 
	-- signal N2_30_52 : std_logic;
	-- signal N2_31_53 : std_logic;
	FA136 : full_adder port map (N0_45_52,N0_46_52,N0_47_52,N2_30_52,N2_31_53);
-- In matrix 1 adding HA to column 52 
	-- signal N2_32_52 : std_logic;
	-- signal N2_33_53 : std_logic;
	HA17 : half_adder port map (N0_48_52,N0_49_52,N2_32_52,N2_33_53);
-- In matrix 1 adding FA to column 53 
	-- signal N2_0_53 : std_logic;
	-- signal N2_1_54 : std_logic;
	FA137 : full_adder port map (N0_1_53,N0_2_53,N0_3_53,N2_0_53,N2_1_54);
-- In matrix 1 adding FA to column 53 
	-- signal N2_2_53 : std_logic;
	-- signal N2_3_54 : std_logic;
	FA138 : full_adder port map (N0_4_53,N0_5_53,N0_6_53,N2_2_53,N2_3_54);
-- In matrix 1 adding FA to column 53 
	-- signal N2_4_53 : std_logic;
	-- signal N2_5_54 : std_logic;
	FA139 : full_adder port map (N0_7_53,N0_8_53,N0_9_53,N2_4_53,N2_5_54);
-- In matrix 1 adding FA to column 53 
	-- signal N2_6_53 : std_logic;
	-- signal N2_7_54 : std_logic;
	FA140 : full_adder port map (N0_10_53,N0_11_53,N0_12_53,N2_6_53,N2_7_54);
-- In matrix 1 adding FA to column 53 
	-- signal N2_8_53 : std_logic;
	-- signal N2_9_54 : std_logic;
	FA141 : full_adder port map (N0_13_53,N0_14_53,N0_15_53,N2_8_53,N2_9_54);
-- In matrix 1 adding FA to column 53 
	-- signal N2_10_53 : std_logic;
	-- signal N2_11_54 : std_logic;
	FA142 : full_adder port map (N0_16_53,N0_17_53,N0_18_53,N2_10_53,N2_11_54);
-- In matrix 1 adding FA to column 53 
	-- signal N2_12_53 : std_logic;
	-- signal N2_13_54 : std_logic;
	FA143 : full_adder port map (N0_19_53,N0_20_53,N0_21_53,N2_12_53,N2_13_54);
-- In matrix 1 adding FA to column 53 
	-- signal N2_14_53 : std_logic;
	-- signal N2_15_54 : std_logic;
	FA144 : full_adder port map (N0_22_53,N0_23_53,N0_24_53,N2_14_53,N2_15_54);
-- In matrix 1 adding FA to column 53 
	-- signal N2_16_53 : std_logic;
	-- signal N2_17_54 : std_logic;
	FA145 : full_adder port map (N0_25_53,N0_26_53,N0_27_53,N2_16_53,N2_17_54);
-- In matrix 1 adding FA to column 53 
	-- signal N2_18_53 : std_logic;
	-- signal N2_19_54 : std_logic;
	FA146 : full_adder port map (N0_28_53,N0_29_53,N0_30_53,N2_18_53,N2_19_54);
-- In matrix 1 adding FA to column 53 
	-- signal N2_20_53 : std_logic;
	-- signal N2_21_54 : std_logic;
	FA147 : full_adder port map (N0_31_53,N0_32_53,N0_33_53,N2_20_53,N2_21_54);
-- In matrix 1 adding FA to column 53 
	-- signal N2_22_53 : std_logic;
	-- signal N2_23_54 : std_logic;
	FA148 : full_adder port map (N0_34_53,N0_35_53,N0_36_53,N2_22_53,N2_23_54);
-- In matrix 1 adding FA to column 53 
	-- signal N2_24_53 : std_logic;
	-- signal N2_25_54 : std_logic;
	FA149 : full_adder port map (N0_37_53,N0_38_53,N0_39_53,N2_24_53,N2_25_54);
-- In matrix 1 adding FA to column 53 
	-- signal N2_26_53 : std_logic;
	-- signal N2_27_54 : std_logic;
	FA150 : full_adder port map (N0_40_53,N0_41_53,N0_42_53,N2_26_53,N2_27_54);
-- In matrix 1 adding FA to column 53 
	-- signal N2_28_53 : std_logic;
	-- signal N2_29_54 : std_logic;
	FA151 : full_adder port map (N0_43_53,N0_44_53,N0_45_53,N2_28_53,N2_29_54);
-- In matrix 1 adding FA to column 53 
	-- signal N2_30_53 : std_logic;
	-- signal N2_31_54 : std_logic;
	FA152 : full_adder port map (N0_46_53,N0_47_53,N0_48_53,N2_30_53,N2_31_54);
-- In matrix 1 adding HA to column 53 
	-- signal N2_32_53 : std_logic;
	-- signal N2_33_54 : std_logic;
	HA18 : half_adder port map (N0_49_53,N0_50_53,N2_32_53,N2_33_54);
-- In matrix 1 adding FA to column 54 
	-- signal N2_0_54 : std_logic;
	-- signal N2_1_55 : std_logic;
	FA153 : full_adder port map (N0_2_54,N0_3_54,N0_4_54,N2_0_54,N2_1_55);
-- In matrix 1 adding FA to column 54 
	-- signal N2_2_54 : std_logic;
	-- signal N2_3_55 : std_logic;
	FA154 : full_adder port map (N0_5_54,N0_6_54,N0_7_54,N2_2_54,N2_3_55);
-- In matrix 1 adding FA to column 54 
	-- signal N2_4_54 : std_logic;
	-- signal N2_5_55 : std_logic;
	FA155 : full_adder port map (N0_8_54,N0_9_54,N0_10_54,N2_4_54,N2_5_55);
-- In matrix 1 adding FA to column 54 
	-- signal N2_6_54 : std_logic;
	-- signal N2_7_55 : std_logic;
	FA156 : full_adder port map (N0_11_54,N0_12_54,N0_13_54,N2_6_54,N2_7_55);
-- In matrix 1 adding FA to column 54 
	-- signal N2_8_54 : std_logic;
	-- signal N2_9_55 : std_logic;
	FA157 : full_adder port map (N0_14_54,N0_15_54,N0_16_54,N2_8_54,N2_9_55);
-- In matrix 1 adding FA to column 54 
	-- signal N2_10_54 : std_logic;
	-- signal N2_11_55 : std_logic;
	FA158 : full_adder port map (N0_17_54,N0_18_54,N0_19_54,N2_10_54,N2_11_55);
-- In matrix 1 adding FA to column 54 
	-- signal N2_12_54 : std_logic;
	-- signal N2_13_55 : std_logic;
	FA159 : full_adder port map (N0_20_54,N0_21_54,N0_22_54,N2_12_54,N2_13_55);
-- In matrix 1 adding FA to column 54 
	-- signal N2_14_54 : std_logic;
	-- signal N2_15_55 : std_logic;
	FA160 : full_adder port map (N0_23_54,N0_24_54,N0_25_54,N2_14_54,N2_15_55);
-- In matrix 1 adding FA to column 54 
	-- signal N2_16_54 : std_logic;
	-- signal N2_17_55 : std_logic;
	FA161 : full_adder port map (N0_26_54,N0_27_54,N0_28_54,N2_16_54,N2_17_55);
-- In matrix 1 adding FA to column 54 
	-- signal N2_18_54 : std_logic;
	-- signal N2_19_55 : std_logic;
	FA162 : full_adder port map (N0_29_54,N0_30_54,N0_31_54,N2_18_54,N2_19_55);
-- In matrix 1 adding FA to column 54 
	-- signal N2_20_54 : std_logic;
	-- signal N2_21_55 : std_logic;
	FA163 : full_adder port map (N0_32_54,N0_33_54,N0_34_54,N2_20_54,N2_21_55);
-- In matrix 1 adding FA to column 54 
	-- signal N2_22_54 : std_logic;
	-- signal N2_23_55 : std_logic;
	FA164 : full_adder port map (N0_35_54,N0_36_54,N0_37_54,N2_22_54,N2_23_55);
-- In matrix 1 adding FA to column 54 
	-- signal N2_24_54 : std_logic;
	-- signal N2_25_55 : std_logic;
	FA165 : full_adder port map (N0_38_54,N0_39_54,N0_40_54,N2_24_54,N2_25_55);
-- In matrix 1 adding FA to column 54 
	-- signal N2_26_54 : std_logic;
	-- signal N2_27_55 : std_logic;
	FA166 : full_adder port map (N0_41_54,N0_42_54,N0_43_54,N2_26_54,N2_27_55);
-- In matrix 1 adding FA to column 54 
	-- signal N2_28_54 : std_logic;
	-- signal N2_29_55 : std_logic;
	FA167 : full_adder port map (N0_44_54,N0_45_54,N0_46_54,N2_28_54,N2_29_55);
-- In matrix 1 adding FA to column 54 
	-- signal N2_30_54 : std_logic;
	-- signal N2_31_55 : std_logic;
	FA168 : full_adder port map (N0_47_54,N0_48_54,N0_49_54,N2_30_54,N2_31_55);
-- In matrix 1 adding FA to column 55 
	-- signal N2_0_55 : std_logic;
	-- signal N2_1_56 : std_logic;
	FA169 : full_adder port map (N0_3_55,N0_4_55,N0_5_55,N2_0_55,N2_1_56);
-- In matrix 1 adding FA to column 55 
	-- signal N2_2_55 : std_logic;
	-- signal N2_3_56 : std_logic;
	FA170 : full_adder port map (N0_6_55,N0_7_55,N0_8_55,N2_2_55,N2_3_56);
-- In matrix 1 adding FA to column 55 
	-- signal N2_4_55 : std_logic;
	-- signal N2_5_56 : std_logic;
	FA171 : full_adder port map (N0_9_55,N0_10_55,N0_11_55,N2_4_55,N2_5_56);
-- In matrix 1 adding FA to column 55 
	-- signal N2_6_55 : std_logic;
	-- signal N2_7_56 : std_logic;
	FA172 : full_adder port map (N0_12_55,N0_13_55,N0_14_55,N2_6_55,N2_7_56);
-- In matrix 1 adding FA to column 55 
	-- signal N2_8_55 : std_logic;
	-- signal N2_9_56 : std_logic;
	FA173 : full_adder port map (N0_15_55,N0_16_55,N0_17_55,N2_8_55,N2_9_56);
-- In matrix 1 adding FA to column 55 
	-- signal N2_10_55 : std_logic;
	-- signal N2_11_56 : std_logic;
	FA174 : full_adder port map (N0_18_55,N0_19_55,N0_20_55,N2_10_55,N2_11_56);
-- In matrix 1 adding FA to column 55 
	-- signal N2_12_55 : std_logic;
	-- signal N2_13_56 : std_logic;
	FA175 : full_adder port map (N0_21_55,N0_22_55,N0_23_55,N2_12_55,N2_13_56);
-- In matrix 1 adding FA to column 55 
	-- signal N2_14_55 : std_logic;
	-- signal N2_15_56 : std_logic;
	FA176 : full_adder port map (N0_24_55,N0_25_55,N0_26_55,N2_14_55,N2_15_56);
-- In matrix 1 adding FA to column 55 
	-- signal N2_16_55 : std_logic;
	-- signal N2_17_56 : std_logic;
	FA177 : full_adder port map (N0_27_55,N0_28_55,N0_29_55,N2_16_55,N2_17_56);
-- In matrix 1 adding FA to column 55 
	-- signal N2_18_55 : std_logic;
	-- signal N2_19_56 : std_logic;
	FA178 : full_adder port map (N0_30_55,N0_31_55,N0_32_55,N2_18_55,N2_19_56);
-- In matrix 1 adding FA to column 55 
	-- signal N2_20_55 : std_logic;
	-- signal N2_21_56 : std_logic;
	FA179 : full_adder port map (N0_33_55,N0_34_55,N0_35_55,N2_20_55,N2_21_56);
-- In matrix 1 adding FA to column 55 
	-- signal N2_22_55 : std_logic;
	-- signal N2_23_56 : std_logic;
	FA180 : full_adder port map (N0_36_55,N0_37_55,N0_38_55,N2_22_55,N2_23_56);
-- In matrix 1 adding FA to column 55 
	-- signal N2_24_55 : std_logic;
	-- signal N2_25_56 : std_logic;
	FA181 : full_adder port map (N0_39_55,N0_40_55,N0_41_55,N2_24_55,N2_25_56);
-- In matrix 1 adding FA to column 55 
	-- signal N2_26_55 : std_logic;
	-- signal N2_27_56 : std_logic;
	FA182 : full_adder port map (N0_42_55,N0_43_55,N0_44_55,N2_26_55,N2_27_56);
-- In matrix 1 adding FA to column 55 
	-- signal N2_28_55 : std_logic;
	-- signal N2_29_56 : std_logic;
	FA183 : full_adder port map (N0_45_55,N0_46_55,N0_47_55,N2_28_55,N2_29_56);
-- In matrix 1 adding FA to column 56 
	-- signal N2_0_56 : std_logic;
	-- signal N2_1_57 : std_logic;
	FA184 : full_adder port map (N0_4_56,N0_5_56,N0_6_56,N2_0_56,N2_1_57);
-- In matrix 1 adding FA to column 56 
	-- signal N2_2_56 : std_logic;
	-- signal N2_3_57 : std_logic;
	FA185 : full_adder port map (N0_7_56,N0_8_56,N0_9_56,N2_2_56,N2_3_57);
-- In matrix 1 adding FA to column 56 
	-- signal N2_4_56 : std_logic;
	-- signal N2_5_57 : std_logic;
	FA186 : full_adder port map (N0_10_56,N0_11_56,N0_12_56,N2_4_56,N2_5_57);
-- In matrix 1 adding FA to column 56 
	-- signal N2_6_56 : std_logic;
	-- signal N2_7_57 : std_logic;
	FA187 : full_adder port map (N0_13_56,N0_14_56,N0_15_56,N2_6_56,N2_7_57);
-- In matrix 1 adding FA to column 56 
	-- signal N2_8_56 : std_logic;
	-- signal N2_9_57 : std_logic;
	FA188 : full_adder port map (N0_16_56,N0_17_56,N0_18_56,N2_8_56,N2_9_57);
-- In matrix 1 adding FA to column 56 
	-- signal N2_10_56 : std_logic;
	-- signal N2_11_57 : std_logic;
	FA189 : full_adder port map (N0_19_56,N0_20_56,N0_21_56,N2_10_56,N2_11_57);
-- In matrix 1 adding FA to column 56 
	-- signal N2_12_56 : std_logic;
	-- signal N2_13_57 : std_logic;
	FA190 : full_adder port map (N0_22_56,N0_23_56,N0_24_56,N2_12_56,N2_13_57);
-- In matrix 1 adding FA to column 56 
	-- signal N2_14_56 : std_logic;
	-- signal N2_15_57 : std_logic;
	FA191 : full_adder port map (N0_25_56,N0_26_56,N0_27_56,N2_14_56,N2_15_57);
-- In matrix 1 adding FA to column 56 
	-- signal N2_16_56 : std_logic;
	-- signal N2_17_57 : std_logic;
	FA192 : full_adder port map (N0_28_56,N0_29_56,N0_30_56,N2_16_56,N2_17_57);
-- In matrix 1 adding FA to column 56 
	-- signal N2_18_56 : std_logic;
	-- signal N2_19_57 : std_logic;
	FA193 : full_adder port map (N0_31_56,N0_32_56,N0_33_56,N2_18_56,N2_19_57);
-- In matrix 1 adding FA to column 56 
	-- signal N2_20_56 : std_logic;
	-- signal N2_21_57 : std_logic;
	FA194 : full_adder port map (N0_34_56,N0_35_56,N0_36_56,N2_20_56,N2_21_57);
-- In matrix 1 adding FA to column 56 
	-- signal N2_22_56 : std_logic;
	-- signal N2_23_57 : std_logic;
	FA195 : full_adder port map (N0_37_56,N0_38_56,N0_39_56,N2_22_56,N2_23_57);
-- In matrix 1 adding FA to column 56 
	-- signal N2_24_56 : std_logic;
	-- signal N2_25_57 : std_logic;
	FA196 : full_adder port map (N0_40_56,N0_41_56,N0_42_56,N2_24_56,N2_25_57);
-- In matrix 1 adding FA to column 56 
	-- signal N2_26_56 : std_logic;
	-- signal N2_27_57 : std_logic;
	FA197 : full_adder port map (N0_43_56,N0_44_56,N0_45_56,N2_26_56,N2_27_57);
-- In matrix 1 adding FA to column 57 
	-- signal N2_0_57 : std_logic;
	-- signal N2_1_58 : std_logic;
	FA198 : full_adder port map (N0_5_57,N0_6_57,N0_7_57,N2_0_57,N2_1_58);
-- In matrix 1 adding FA to column 57 
	-- signal N2_2_57 : std_logic;
	-- signal N2_3_58 : std_logic;
	FA199 : full_adder port map (N0_8_57,N0_9_57,N0_10_57,N2_2_57,N2_3_58);
-- In matrix 1 adding FA to column 57 
	-- signal N2_4_57 : std_logic;
	-- signal N2_5_58 : std_logic;
	FA200 : full_adder port map (N0_11_57,N0_12_57,N0_13_57,N2_4_57,N2_5_58);
-- In matrix 1 adding FA to column 57 
	-- signal N2_6_57 : std_logic;
	-- signal N2_7_58 : std_logic;
	FA201 : full_adder port map (N0_14_57,N0_15_57,N0_16_57,N2_6_57,N2_7_58);
-- In matrix 1 adding FA to column 57 
	-- signal N2_8_57 : std_logic;
	-- signal N2_9_58 : std_logic;
	FA202 : full_adder port map (N0_17_57,N0_18_57,N0_19_57,N2_8_57,N2_9_58);
-- In matrix 1 adding FA to column 57 
	-- signal N2_10_57 : std_logic;
	-- signal N2_11_58 : std_logic;
	FA203 : full_adder port map (N0_20_57,N0_21_57,N0_22_57,N2_10_57,N2_11_58);
-- In matrix 1 adding FA to column 57 
	-- signal N2_12_57 : std_logic;
	-- signal N2_13_58 : std_logic;
	FA204 : full_adder port map (N0_23_57,N0_24_57,N0_25_57,N2_12_57,N2_13_58);
-- In matrix 1 adding FA to column 57 
	-- signal N2_14_57 : std_logic;
	-- signal N2_15_58 : std_logic;
	FA205 : full_adder port map (N0_26_57,N0_27_57,N0_28_57,N2_14_57,N2_15_58);
-- In matrix 1 adding FA to column 57 
	-- signal N2_16_57 : std_logic;
	-- signal N2_17_58 : std_logic;
	FA206 : full_adder port map (N0_29_57,N0_30_57,N0_31_57,N2_16_57,N2_17_58);
-- In matrix 1 adding FA to column 57 
	-- signal N2_18_57 : std_logic;
	-- signal N2_19_58 : std_logic;
	FA207 : full_adder port map (N0_32_57,N0_33_57,N0_34_57,N2_18_57,N2_19_58);
-- In matrix 1 adding FA to column 57 
	-- signal N2_20_57 : std_logic;
	-- signal N2_21_58 : std_logic;
	FA208 : full_adder port map (N0_35_57,N0_36_57,N0_37_57,N2_20_57,N2_21_58);
-- In matrix 1 adding FA to column 57 
	-- signal N2_22_57 : std_logic;
	-- signal N2_23_58 : std_logic;
	FA209 : full_adder port map (N0_38_57,N0_39_57,N0_40_57,N2_22_57,N2_23_58);
-- In matrix 1 adding FA to column 57 
	-- signal N2_24_57 : std_logic;
	-- signal N2_25_58 : std_logic;
	FA210 : full_adder port map (N0_41_57,N0_42_57,N0_43_57,N2_24_57,N2_25_58);
-- In matrix 1 adding FA to column 58 
	-- signal N2_0_58 : std_logic;
	-- signal N2_1_59 : std_logic;
	FA211 : full_adder port map (N0_6_58,N0_7_58,N0_8_58,N2_0_58,N2_1_59);
-- In matrix 1 adding FA to column 58 
	-- signal N2_2_58 : std_logic;
	-- signal N2_3_59 : std_logic;
	FA212 : full_adder port map (N0_9_58,N0_10_58,N0_11_58,N2_2_58,N2_3_59);
-- In matrix 1 adding FA to column 58 
	-- signal N2_4_58 : std_logic;
	-- signal N2_5_59 : std_logic;
	FA213 : full_adder port map (N0_12_58,N0_13_58,N0_14_58,N2_4_58,N2_5_59);
-- In matrix 1 adding FA to column 58 
	-- signal N2_6_58 : std_logic;
	-- signal N2_7_59 : std_logic;
	FA214 : full_adder port map (N0_15_58,N0_16_58,N0_17_58,N2_6_58,N2_7_59);
-- In matrix 1 adding FA to column 58 
	-- signal N2_8_58 : std_logic;
	-- signal N2_9_59 : std_logic;
	FA215 : full_adder port map (N0_18_58,N0_19_58,N0_20_58,N2_8_58,N2_9_59);
-- In matrix 1 adding FA to column 58 
	-- signal N2_10_58 : std_logic;
	-- signal N2_11_59 : std_logic;
	FA216 : full_adder port map (N0_21_58,N0_22_58,N0_23_58,N2_10_58,N2_11_59);
-- In matrix 1 adding FA to column 58 
	-- signal N2_12_58 : std_logic;
	-- signal N2_13_59 : std_logic;
	FA217 : full_adder port map (N0_24_58,N0_25_58,N0_26_58,N2_12_58,N2_13_59);
-- In matrix 1 adding FA to column 58 
	-- signal N2_14_58 : std_logic;
	-- signal N2_15_59 : std_logic;
	FA218 : full_adder port map (N0_27_58,N0_28_58,N0_29_58,N2_14_58,N2_15_59);
-- In matrix 1 adding FA to column 58 
	-- signal N2_16_58 : std_logic;
	-- signal N2_17_59 : std_logic;
	FA219 : full_adder port map (N0_30_58,N0_31_58,N0_32_58,N2_16_58,N2_17_59);
-- In matrix 1 adding FA to column 58 
	-- signal N2_18_58 : std_logic;
	-- signal N2_19_59 : std_logic;
	FA220 : full_adder port map (N0_33_58,N0_34_58,N0_35_58,N2_18_58,N2_19_59);
-- In matrix 1 adding FA to column 58 
	-- signal N2_20_58 : std_logic;
	-- signal N2_21_59 : std_logic;
	FA221 : full_adder port map (N0_36_58,N0_37_58,N0_38_58,N2_20_58,N2_21_59);
-- In matrix 1 adding FA to column 58 
	-- signal N2_22_58 : std_logic;
	-- signal N2_23_59 : std_logic;
	FA222 : full_adder port map (N0_39_58,N0_40_58,N0_41_58,N2_22_58,N2_23_59);
-- In matrix 1 adding FA to column 59 
	-- signal N2_0_59 : std_logic;
	-- signal N2_1_60 : std_logic;
	FA223 : full_adder port map (N0_7_59,N0_8_59,N0_9_59,N2_0_59,N2_1_60);
-- In matrix 1 adding FA to column 59 
	-- signal N2_2_59 : std_logic;
	-- signal N2_3_60 : std_logic;
	FA224 : full_adder port map (N0_10_59,N0_11_59,N0_12_59,N2_2_59,N2_3_60);
-- In matrix 1 adding FA to column 59 
	-- signal N2_4_59 : std_logic;
	-- signal N2_5_60 : std_logic;
	FA225 : full_adder port map (N0_13_59,N0_14_59,N0_15_59,N2_4_59,N2_5_60);
-- In matrix 1 adding FA to column 59 
	-- signal N2_6_59 : std_logic;
	-- signal N2_7_60 : std_logic;
	FA226 : full_adder port map (N0_16_59,N0_17_59,N0_18_59,N2_6_59,N2_7_60);
-- In matrix 1 adding FA to column 59 
	-- signal N2_8_59 : std_logic;
	-- signal N2_9_60 : std_logic;
	FA227 : full_adder port map (N0_19_59,N0_20_59,N0_21_59,N2_8_59,N2_9_60);
-- In matrix 1 adding FA to column 59 
	-- signal N2_10_59 : std_logic;
	-- signal N2_11_60 : std_logic;
	FA228 : full_adder port map (N0_22_59,N0_23_59,N0_24_59,N2_10_59,N2_11_60);
-- In matrix 1 adding FA to column 59 
	-- signal N2_12_59 : std_logic;
	-- signal N2_13_60 : std_logic;
	FA229 : full_adder port map (N0_25_59,N0_26_59,N0_27_59,N2_12_59,N2_13_60);
-- In matrix 1 adding FA to column 59 
	-- signal N2_14_59 : std_logic;
	-- signal N2_15_60 : std_logic;
	FA230 : full_adder port map (N0_28_59,N0_29_59,N0_30_59,N2_14_59,N2_15_60);
-- In matrix 1 adding FA to column 59 
	-- signal N2_16_59 : std_logic;
	-- signal N2_17_60 : std_logic;
	FA231 : full_adder port map (N0_31_59,N0_32_59,N0_33_59,N2_16_59,N2_17_60);
-- In matrix 1 adding FA to column 59 
	-- signal N2_18_59 : std_logic;
	-- signal N2_19_60 : std_logic;
	FA232 : full_adder port map (N0_34_59,N0_35_59,N0_36_59,N2_18_59,N2_19_60);
-- In matrix 1 adding FA to column 59 
	-- signal N2_20_59 : std_logic;
	-- signal N2_21_60 : std_logic;
	FA233 : full_adder port map (N0_37_59,N0_38_59,N0_39_59,N2_20_59,N2_21_60);
-- In matrix 1 adding FA to column 60 
	-- signal N2_0_60 : std_logic;
	-- signal N2_1_61 : std_logic;
	FA234 : full_adder port map (N0_8_60,N0_9_60,N0_10_60,N2_0_60,N2_1_61);
-- In matrix 1 adding FA to column 60 
	-- signal N2_2_60 : std_logic;
	-- signal N2_3_61 : std_logic;
	FA235 : full_adder port map (N0_11_60,N0_12_60,N0_13_60,N2_2_60,N2_3_61);
-- In matrix 1 adding FA to column 60 
	-- signal N2_4_60 : std_logic;
	-- signal N2_5_61 : std_logic;
	FA236 : full_adder port map (N0_14_60,N0_15_60,N0_16_60,N2_4_60,N2_5_61);
-- In matrix 1 adding FA to column 60 
	-- signal N2_6_60 : std_logic;
	-- signal N2_7_61 : std_logic;
	FA237 : full_adder port map (N0_17_60,N0_18_60,N0_19_60,N2_6_60,N2_7_61);
-- In matrix 1 adding FA to column 60 
	-- signal N2_8_60 : std_logic;
	-- signal N2_9_61 : std_logic;
	FA238 : full_adder port map (N0_20_60,N0_21_60,N0_22_60,N2_8_60,N2_9_61);
-- In matrix 1 adding FA to column 60 
	-- signal N2_10_60 : std_logic;
	-- signal N2_11_61 : std_logic;
	FA239 : full_adder port map (N0_23_60,N0_24_60,N0_25_60,N2_10_60,N2_11_61);
-- In matrix 1 adding FA to column 60 
	-- signal N2_12_60 : std_logic;
	-- signal N2_13_61 : std_logic;
	FA240 : full_adder port map (N0_26_60,N0_27_60,N0_28_60,N2_12_60,N2_13_61);
-- In matrix 1 adding FA to column 60 
	-- signal N2_14_60 : std_logic;
	-- signal N2_15_61 : std_logic;
	FA241 : full_adder port map (N0_29_60,N0_30_60,N0_31_60,N2_14_60,N2_15_61);
-- In matrix 1 adding FA to column 60 
	-- signal N2_16_60 : std_logic;
	-- signal N2_17_61 : std_logic;
	FA242 : full_adder port map (N0_32_60,N0_33_60,N0_34_60,N2_16_60,N2_17_61);
-- In matrix 1 adding FA to column 60 
	-- signal N2_18_60 : std_logic;
	-- signal N2_19_61 : std_logic;
	FA243 : full_adder port map (N0_35_60,N0_36_60,N0_37_60,N2_18_60,N2_19_61);
-- In matrix 1 adding FA to column 61 
	-- signal N2_0_61 : std_logic;
	-- signal N2_1_62 : std_logic;
	FA244 : full_adder port map (N0_9_61,N0_10_61,N0_11_61,N2_0_61,N2_1_62);
-- In matrix 1 adding FA to column 61 
	-- signal N2_2_61 : std_logic;
	-- signal N2_3_62 : std_logic;
	FA245 : full_adder port map (N0_12_61,N0_13_61,N0_14_61,N2_2_61,N2_3_62);
-- In matrix 1 adding FA to column 61 
	-- signal N2_4_61 : std_logic;
	-- signal N2_5_62 : std_logic;
	FA246 : full_adder port map (N0_15_61,N0_16_61,N0_17_61,N2_4_61,N2_5_62);
-- In matrix 1 adding FA to column 61 
	-- signal N2_6_61 : std_logic;
	-- signal N2_7_62 : std_logic;
	FA247 : full_adder port map (N0_18_61,N0_19_61,N0_20_61,N2_6_61,N2_7_62);
-- In matrix 1 adding FA to column 61 
	-- signal N2_8_61 : std_logic;
	-- signal N2_9_62 : std_logic;
	FA248 : full_adder port map (N0_21_61,N0_22_61,N0_23_61,N2_8_61,N2_9_62);
-- In matrix 1 adding FA to column 61 
	-- signal N2_10_61 : std_logic;
	-- signal N2_11_62 : std_logic;
	FA249 : full_adder port map (N0_24_61,N0_25_61,N0_26_61,N2_10_61,N2_11_62);
-- In matrix 1 adding FA to column 61 
	-- signal N2_12_61 : std_logic;
	-- signal N2_13_62 : std_logic;
	FA250 : full_adder port map (N0_27_61,N0_28_61,N0_29_61,N2_12_61,N2_13_62);
-- In matrix 1 adding FA to column 61 
	-- signal N2_14_61 : std_logic;
	-- signal N2_15_62 : std_logic;
	FA251 : full_adder port map (N0_30_61,N0_31_61,N0_32_61,N2_14_61,N2_15_62);
-- In matrix 1 adding FA to column 61 
	-- signal N2_16_61 : std_logic;
	-- signal N2_17_62 : std_logic;
	FA252 : full_adder port map (N0_33_61,N0_34_61,N0_35_61,N2_16_61,N2_17_62);
-- In matrix 1 adding FA to column 62 
	-- signal N2_0_62 : std_logic;
	-- signal N2_1_63 : std_logic;
	FA253 : full_adder port map (N0_10_62,N0_11_62,N0_12_62,N2_0_62,N2_1_63);
-- In matrix 1 adding FA to column 62 
	-- signal N2_2_62 : std_logic;
	-- signal N2_3_63 : std_logic;
	FA254 : full_adder port map (N0_13_62,N0_14_62,N0_15_62,N2_2_62,N2_3_63);
-- In matrix 1 adding FA to column 62 
	-- signal N2_4_62 : std_logic;
	-- signal N2_5_63 : std_logic;
	FA255 : full_adder port map (N0_16_62,N0_17_62,N0_18_62,N2_4_62,N2_5_63);
-- In matrix 1 adding FA to column 62 
	-- signal N2_6_62 : std_logic;
	-- signal N2_7_63 : std_logic;
	FA256 : full_adder port map (N0_19_62,N0_20_62,N0_21_62,N2_6_62,N2_7_63);
-- In matrix 1 adding FA to column 62 
	-- signal N2_8_62 : std_logic;
	-- signal N2_9_63 : std_logic;
	FA257 : full_adder port map (N0_22_62,N0_23_62,N0_24_62,N2_8_62,N2_9_63);
-- In matrix 1 adding FA to column 62 
	-- signal N2_10_62 : std_logic;
	-- signal N2_11_63 : std_logic;
	FA258 : full_adder port map (N0_25_62,N0_26_62,N0_27_62,N2_10_62,N2_11_63);
-- In matrix 1 adding FA to column 62 
	-- signal N2_12_62 : std_logic;
	-- signal N2_13_63 : std_logic;
	FA259 : full_adder port map (N0_28_62,N0_29_62,N0_30_62,N2_12_62,N2_13_63);
-- In matrix 1 adding FA to column 62 
	-- signal N2_14_62 : std_logic;
	-- signal N2_15_63 : std_logic;
	FA260 : full_adder port map (N0_31_62,N0_32_62,N0_33_62,N2_14_62,N2_15_63);
-- In matrix 1 adding FA to column 63 
	-- signal N2_0_63 : std_logic;
	-- signal N2_1_64 : std_logic;
	FA261 : full_adder port map (N0_11_63,N0_12_63,N0_13_63,N2_0_63,N2_1_64);
-- In matrix 1 adding FA to column 63 
	-- signal N2_2_63 : std_logic;
	-- signal N2_3_64 : std_logic;
	FA262 : full_adder port map (N0_14_63,N0_15_63,N0_16_63,N2_2_63,N2_3_64);
-- In matrix 1 adding FA to column 63 
	-- signal N2_4_63 : std_logic;
	-- signal N2_5_64 : std_logic;
	FA263 : full_adder port map (N0_17_63,N0_18_63,N0_19_63,N2_4_63,N2_5_64);
-- In matrix 1 adding FA to column 63 
	-- signal N2_6_63 : std_logic;
	-- signal N2_7_64 : std_logic;
	FA264 : full_adder port map (N0_20_63,N0_21_63,N0_22_63,N2_6_63,N2_7_64);
-- In matrix 1 adding FA to column 63 
	-- signal N2_8_63 : std_logic;
	-- signal N2_9_64 : std_logic;
	FA265 : full_adder port map (N0_23_63,N0_24_63,N0_25_63,N2_8_63,N2_9_64);
-- In matrix 1 adding FA to column 63 
	-- signal N2_10_63 : std_logic;
	-- signal N2_11_64 : std_logic;
	FA266 : full_adder port map (N0_26_63,N0_27_63,N0_28_63,N2_10_63,N2_11_64);
-- In matrix 1 adding FA to column 63 
	-- signal N2_12_63 : std_logic;
	-- signal N2_13_64 : std_logic;
	FA267 : full_adder port map (N0_29_63,N0_30_63,N0_31_63,N2_12_63,N2_13_64);
-- In matrix 1 adding FA to column 64 
	-- signal N2_0_64 : std_logic;
	-- signal N2_1_65 : std_logic;
	FA268 : full_adder port map (N0_12_64,N0_13_64,N0_14_64,N2_0_64,N2_1_65);
-- In matrix 1 adding FA to column 64 
	-- signal N2_2_64 : std_logic;
	-- signal N2_3_65 : std_logic;
	FA269 : full_adder port map (N0_15_64,N0_16_64,N0_17_64,N2_2_64,N2_3_65);
-- In matrix 1 adding FA to column 64 
	-- signal N2_4_64 : std_logic;
	-- signal N2_5_65 : std_logic;
	FA270 : full_adder port map (N0_18_64,N0_19_64,N0_20_64,N2_4_64,N2_5_65);
-- In matrix 1 adding FA to column 64 
	-- signal N2_6_64 : std_logic;
	-- signal N2_7_65 : std_logic;
	FA271 : full_adder port map (N0_21_64,N0_22_64,N0_23_64,N2_6_64,N2_7_65);
-- In matrix 1 adding FA to column 64 
	-- signal N2_8_64 : std_logic;
	-- signal N2_9_65 : std_logic;
	FA272 : full_adder port map (N0_24_64,N0_25_64,N0_26_64,N2_8_64,N2_9_65);
-- In matrix 1 adding FA to column 64 
	-- signal N2_10_64 : std_logic;
	-- signal N2_11_65 : std_logic;
	FA273 : full_adder port map (N0_27_64,N0_28_64,N0_29_64,N2_10_64,N2_11_65);
-- In matrix 1 adding FA to column 65 
	-- signal N2_0_65 : std_logic;
	-- signal N2_1_66 : std_logic;
	FA274 : full_adder port map (N0_13_65,N0_14_65,N0_15_65,N2_0_65,N2_1_66);
-- In matrix 1 adding FA to column 65 
	-- signal N2_2_65 : std_logic;
	-- signal N2_3_66 : std_logic;
	FA275 : full_adder port map (N0_16_65,N0_17_65,N0_18_65,N2_2_65,N2_3_66);
-- In matrix 1 adding FA to column 65 
	-- signal N2_4_65 : std_logic;
	-- signal N2_5_66 : std_logic;
	FA276 : full_adder port map (N0_19_65,N0_20_65,N0_21_65,N2_4_65,N2_5_66);
-- In matrix 1 adding FA to column 65 
	-- signal N2_6_65 : std_logic;
	-- signal N2_7_66 : std_logic;
	FA277 : full_adder port map (N0_22_65,N0_23_65,N0_24_65,N2_6_65,N2_7_66);
-- In matrix 1 adding FA to column 65 
	-- signal N2_8_65 : std_logic;
	-- signal N2_9_66 : std_logic;
	FA278 : full_adder port map (N0_25_65,N0_26_65,N0_27_65,N2_8_65,N2_9_66);
-- In matrix 1 adding FA to column 66 
	-- signal N2_0_66 : std_logic;
	-- signal N2_1_67 : std_logic;
	FA279 : full_adder port map (N0_14_66,N0_15_66,N0_16_66,N2_0_66,N2_1_67);
-- In matrix 1 adding FA to column 66 
	-- signal N2_2_66 : std_logic;
	-- signal N2_3_67 : std_logic;
	FA280 : full_adder port map (N0_17_66,N0_18_66,N0_19_66,N2_2_66,N2_3_67);
-- In matrix 1 adding FA to column 66 
	-- signal N2_4_66 : std_logic;
	-- signal N2_5_67 : std_logic;
	FA281 : full_adder port map (N0_20_66,N0_21_66,N0_22_66,N2_4_66,N2_5_67);
-- In matrix 1 adding FA to column 66 
	-- signal N2_6_66 : std_logic;
	-- signal N2_7_67 : std_logic;
	FA282 : full_adder port map (N0_23_66,N0_24_66,N0_25_66,N2_6_66,N2_7_67);
-- In matrix 1 adding FA to column 67 
	-- signal N2_0_67 : std_logic;
	-- signal N2_1_68 : std_logic;
	FA283 : full_adder port map (N0_15_67,N0_16_67,N0_17_67,N2_0_67,N2_1_68);
-- In matrix 1 adding FA to column 67 
	-- signal N2_2_67 : std_logic;
	-- signal N2_3_68 : std_logic;
	FA284 : full_adder port map (N0_18_67,N0_19_67,N0_20_67,N2_2_67,N2_3_68);
-- In matrix 1 adding FA to column 67 
	-- signal N2_4_67 : std_logic;
	-- signal N2_5_68 : std_logic;
	FA285 : full_adder port map (N0_21_67,N0_22_67,N0_23_67,N2_4_67,N2_5_68);
-- In matrix 1 adding FA to column 68 
	-- signal N2_0_68 : std_logic;
	-- signal N2_1_69 : std_logic;
	FA286 : full_adder port map (N0_16_68,N0_17_68,N0_18_68,N2_0_68,N2_1_69);
-- In matrix 1 adding FA to column 68 
	-- signal N2_2_68 : std_logic;
	-- signal N2_3_69 : std_logic;
	FA287 : full_adder port map (N0_19_68,N0_20_68,N0_21_68,N2_2_68,N2_3_69);
-- In matrix 1 adding FA to column 69 
	-- signal N2_0_69 : std_logic;
	-- signal N2_1_70 : std_logic;
	FA288 : full_adder port map (N0_17_69,N0_18_69,N0_19_69,N2_0_69,N2_1_70);
	-- Elements from matrix 2 
-- In matrix 2 adding HA to column 24 
	-- signal N3_0_24 : std_logic;
	-- signal N3_1_25 : std_logic;
	HA19 : half_adder port map (N0_0_24,N0_1_24,N3_0_24,N3_1_25);
-- In matrix 2 adding FA to column 25 
	-- signal N3_0_25 : std_logic;
	-- signal N3_1_26 : std_logic;
	FA289 : full_adder port map (N0_0_25,N0_1_25,N0_2_25,N3_0_25,N3_1_26);
-- In matrix 2 adding HA to column 25 
	-- signal N3_2_25 : std_logic;
	-- signal N3_3_26 : std_logic;
	HA20 : half_adder port map (N0_3_25,N0_4_25,N3_2_25,N3_3_26);
-- In matrix 2 adding FA to column 26 
	-- signal N3_0_26 : std_logic;
	-- signal N3_1_27 : std_logic;
	FA290 : full_adder port map (N0_0_26,N0_1_26,N0_2_26,N3_0_26,N3_1_27);
-- In matrix 2 adding FA to column 26 
	-- signal N3_2_26 : std_logic;
	-- signal N3_3_27 : std_logic;
	FA291 : full_adder port map (N0_3_26,N0_4_26,N0_5_26,N3_2_26,N3_3_27);
-- In matrix 2 adding HA to column 26 
	-- signal N3_4_26 : std_logic;
	-- signal N3_5_27 : std_logic;
	HA21 : half_adder port map (N0_6_26,N0_7_26,N3_4_26,N3_5_27);
-- In matrix 2 adding FA to column 27 
	-- signal N3_0_27 : std_logic;
	-- signal N3_1_28 : std_logic;
	FA292 : full_adder port map (N0_0_27,N0_1_27,N0_2_27,N3_0_27,N3_1_28);
-- In matrix 2 adding FA to column 27 
	-- signal N3_2_27 : std_logic;
	-- signal N3_3_28 : std_logic;
	FA293 : full_adder port map (N0_3_27,N0_4_27,N0_5_27,N3_2_27,N3_3_28);
-- In matrix 2 adding FA to column 27 
	-- signal N3_4_27 : std_logic;
	-- signal N3_5_28 : std_logic;
	FA294 : full_adder port map (N0_6_27,N0_7_27,N0_8_27,N3_4_27,N3_5_28);
-- In matrix 2 adding HA to column 27 
	-- signal N3_6_27 : std_logic;
	-- signal N3_7_28 : std_logic;
	HA22 : half_adder port map (N0_9_27,N0_10_27,N3_6_27,N3_7_28);
-- In matrix 2 adding FA to column 28 
	-- signal N3_0_28 : std_logic;
	-- signal N3_1_29 : std_logic;
	FA295 : full_adder port map (N0_0_28,N0_1_28,N0_2_28,N3_0_28,N3_1_29);
-- In matrix 2 adding FA to column 28 
	-- signal N3_2_28 : std_logic;
	-- signal N3_3_29 : std_logic;
	FA296 : full_adder port map (N0_3_28,N0_4_28,N0_5_28,N3_2_28,N3_3_29);
-- In matrix 2 adding FA to column 28 
	-- signal N3_4_28 : std_logic;
	-- signal N3_5_29 : std_logic;
	FA297 : full_adder port map (N0_6_28,N0_7_28,N0_8_28,N3_4_28,N3_5_29);
-- In matrix 2 adding FA to column 28 
	-- signal N3_6_28 : std_logic;
	-- signal N3_7_29 : std_logic;
	FA298 : full_adder port map (N0_9_28,N0_10_28,N0_11_28,N3_6_28,N3_7_29);
-- In matrix 2 adding HA to column 28 
	-- signal N3_8_28 : std_logic;
	-- signal N3_9_29 : std_logic;
	HA23 : half_adder port map (N0_12_28,N0_13_28,N3_8_28,N3_9_29);
-- In matrix 2 adding FA to column 29 
	-- signal N3_0_29 : std_logic;
	-- signal N3_1_30 : std_logic;
	FA299 : full_adder port map (N0_0_29,N0_1_29,N0_2_29,N3_0_29,N3_1_30);
-- In matrix 2 adding FA to column 29 
	-- signal N3_2_29 : std_logic;
	-- signal N3_3_30 : std_logic;
	FA300 : full_adder port map (N0_3_29,N0_4_29,N0_5_29,N3_2_29,N3_3_30);
-- In matrix 2 adding FA to column 29 
	-- signal N3_4_29 : std_logic;
	-- signal N3_5_30 : std_logic;
	FA301 : full_adder port map (N0_6_29,N0_7_29,N0_8_29,N3_4_29,N3_5_30);
-- In matrix 2 adding FA to column 29 
	-- signal N3_6_29 : std_logic;
	-- signal N3_7_30 : std_logic;
	FA302 : full_adder port map (N0_9_29,N0_10_29,N0_11_29,N3_6_29,N3_7_30);
-- In matrix 2 adding FA to column 29 
	-- signal N3_8_29 : std_logic;
	-- signal N3_9_30 : std_logic;
	FA303 : full_adder port map (N0_12_29,N0_13_29,N0_14_29,N3_8_29,N3_9_30);
-- In matrix 2 adding HA to column 29 
	-- signal N3_10_29 : std_logic;
	-- signal N3_11_30 : std_logic;
	HA24 : half_adder port map (N0_15_29,N0_16_29,N3_10_29,N3_11_30);
-- In matrix 2 adding FA to column 30 
	-- signal N3_0_30 : std_logic;
	-- signal N3_1_31 : std_logic;
	FA304 : full_adder port map (N0_0_30,N0_1_30,N0_2_30,N3_0_30,N3_1_31);
-- In matrix 2 adding FA to column 30 
	-- signal N3_2_30 : std_logic;
	-- signal N3_3_31 : std_logic;
	FA305 : full_adder port map (N0_3_30,N0_4_30,N0_5_30,N3_2_30,N3_3_31);
-- In matrix 2 adding FA to column 30 
	-- signal N3_4_30 : std_logic;
	-- signal N3_5_31 : std_logic;
	FA306 : full_adder port map (N0_6_30,N0_7_30,N0_8_30,N3_4_30,N3_5_31);
-- In matrix 2 adding FA to column 30 
	-- signal N3_6_30 : std_logic;
	-- signal N3_7_31 : std_logic;
	FA307 : full_adder port map (N0_9_30,N0_10_30,N0_11_30,N3_6_30,N3_7_31);
-- In matrix 2 adding FA to column 30 
	-- signal N3_8_30 : std_logic;
	-- signal N3_9_31 : std_logic;
	FA308 : full_adder port map (N0_12_30,N0_13_30,N0_14_30,N3_8_30,N3_9_31);
-- In matrix 2 adding FA to column 30 
	-- signal N3_10_30 : std_logic;
	-- signal N3_11_31 : std_logic;
	FA309 : full_adder port map (N0_15_30,N0_16_30,N0_17_30,N3_10_30,N3_11_31);
-- In matrix 2 adding HA to column 30 
	-- signal N3_12_30 : std_logic;
	-- signal N3_13_31 : std_logic;
	HA25 : half_adder port map (N0_18_30,N0_19_30,N3_12_30,N3_13_31);
-- In matrix 2 adding FA to column 31 
	-- signal N3_0_31 : std_logic;
	-- signal N3_1_32 : std_logic;
	FA310 : full_adder port map (N0_0_31,N0_1_31,N0_2_31,N3_0_31,N3_1_32);
-- In matrix 2 adding FA to column 31 
	-- signal N3_2_31 : std_logic;
	-- signal N3_3_32 : std_logic;
	FA311 : full_adder port map (N0_3_31,N0_4_31,N0_5_31,N3_2_31,N3_3_32);
-- In matrix 2 adding FA to column 31 
	-- signal N3_4_31 : std_logic;
	-- signal N3_5_32 : std_logic;
	FA312 : full_adder port map (N0_6_31,N0_7_31,N0_8_31,N3_4_31,N3_5_32);
-- In matrix 2 adding FA to column 31 
	-- signal N3_6_31 : std_logic;
	-- signal N3_7_32 : std_logic;
	FA313 : full_adder port map (N0_9_31,N0_10_31,N0_11_31,N3_6_31,N3_7_32);
-- In matrix 2 adding FA to column 31 
	-- signal N3_8_31 : std_logic;
	-- signal N3_9_32 : std_logic;
	FA314 : full_adder port map (N0_12_31,N0_13_31,N0_14_31,N3_8_31,N3_9_32);
-- In matrix 2 adding FA to column 31 
	-- signal N3_10_31 : std_logic;
	-- signal N3_11_32 : std_logic;
	FA315 : full_adder port map (N0_15_31,N0_16_31,N0_17_31,N3_10_31,N3_11_32);
-- In matrix 2 adding FA to column 31 
	-- signal N3_12_31 : std_logic;
	-- signal N3_13_32 : std_logic;
	FA316 : full_adder port map (N0_18_31,N0_19_31,N0_20_31,N3_12_31,N3_13_32);
-- In matrix 2 adding HA to column 31 
	-- signal N3_14_31 : std_logic;
	-- signal N3_15_32 : std_logic;
	HA26 : half_adder port map (N0_21_31,N0_22_31,N3_14_31,N3_15_32);
-- In matrix 2 adding FA to column 32 
	-- signal N3_0_32 : std_logic;
	-- signal N3_1_33 : std_logic;
	FA317 : full_adder port map (N0_0_32,N0_1_32,N0_2_32,N3_0_32,N3_1_33);
-- In matrix 2 adding FA to column 32 
	-- signal N3_2_32 : std_logic;
	-- signal N3_3_33 : std_logic;
	FA318 : full_adder port map (N0_3_32,N0_4_32,N0_5_32,N3_2_32,N3_3_33);
-- In matrix 2 adding FA to column 32 
	-- signal N3_4_32 : std_logic;
	-- signal N3_5_33 : std_logic;
	FA319 : full_adder port map (N0_6_32,N0_7_32,N0_8_32,N3_4_32,N3_5_33);
-- In matrix 2 adding FA to column 32 
	-- signal N3_6_32 : std_logic;
	-- signal N3_7_33 : std_logic;
	FA320 : full_adder port map (N0_9_32,N0_10_32,N0_11_32,N3_6_32,N3_7_33);
-- In matrix 2 adding FA to column 32 
	-- signal N3_8_32 : std_logic;
	-- signal N3_9_33 : std_logic;
	FA321 : full_adder port map (N0_12_32,N0_13_32,N0_14_32,N3_8_32,N3_9_33);
-- In matrix 2 adding FA to column 32 
	-- signal N3_10_32 : std_logic;
	-- signal N3_11_33 : std_logic;
	FA322 : full_adder port map (N0_15_32,N0_16_32,N0_17_32,N3_10_32,N3_11_33);
-- In matrix 2 adding FA to column 32 
	-- signal N3_12_32 : std_logic;
	-- signal N3_13_33 : std_logic;
	FA323 : full_adder port map (N0_18_32,N0_19_32,N0_20_32,N3_12_32,N3_13_33);
-- In matrix 2 adding FA to column 32 
	-- signal N3_14_32 : std_logic;
	-- signal N3_15_33 : std_logic;
	FA324 : full_adder port map (N0_21_32,N0_22_32,N0_23_32,N3_14_32,N3_15_33);
-- In matrix 2 adding HA to column 32 
	-- signal N3_16_32 : std_logic;
	-- signal N3_17_33 : std_logic;
	HA27 : half_adder port map (N0_24_32,N0_25_32,N3_16_32,N3_17_33);
-- In matrix 2 adding FA to column 33 
	-- signal N3_0_33 : std_logic;
	-- signal N3_1_34 : std_logic;
	FA325 : full_adder port map (N0_0_33,N0_1_33,N0_2_33,N3_0_33,N3_1_34);
-- In matrix 2 adding FA to column 33 
	-- signal N3_2_33 : std_logic;
	-- signal N3_3_34 : std_logic;
	FA326 : full_adder port map (N0_3_33,N0_4_33,N0_5_33,N3_2_33,N3_3_34);
-- In matrix 2 adding FA to column 33 
	-- signal N3_4_33 : std_logic;
	-- signal N3_5_34 : std_logic;
	FA327 : full_adder port map (N0_6_33,N0_7_33,N0_8_33,N3_4_33,N3_5_34);
-- In matrix 2 adding FA to column 33 
	-- signal N3_6_33 : std_logic;
	-- signal N3_7_34 : std_logic;
	FA328 : full_adder port map (N0_9_33,N0_10_33,N0_11_33,N3_6_33,N3_7_34);
-- In matrix 2 adding FA to column 33 
	-- signal N3_8_33 : std_logic;
	-- signal N3_9_34 : std_logic;
	FA329 : full_adder port map (N0_12_33,N0_13_33,N0_14_33,N3_8_33,N3_9_34);
-- In matrix 2 adding FA to column 33 
	-- signal N3_10_33 : std_logic;
	-- signal N3_11_34 : std_logic;
	FA330 : full_adder port map (N0_15_33,N0_16_33,N0_17_33,N3_10_33,N3_11_34);
-- In matrix 2 adding FA to column 33 
	-- signal N3_12_33 : std_logic;
	-- signal N3_13_34 : std_logic;
	FA331 : full_adder port map (N0_18_33,N0_19_33,N0_20_33,N3_12_33,N3_13_34);
-- In matrix 2 adding FA to column 33 
	-- signal N3_14_33 : std_logic;
	-- signal N3_15_34 : std_logic;
	FA332 : full_adder port map (N0_21_33,N0_22_33,N0_23_33,N3_14_33,N3_15_34);
-- In matrix 2 adding FA to column 33 
	-- signal N3_16_33 : std_logic;
	-- signal N3_17_34 : std_logic;
	FA333 : full_adder port map (N0_24_33,N0_25_33,N0_26_33,N3_16_33,N3_17_34);
-- In matrix 2 adding HA to column 33 
	-- signal N3_18_33 : std_logic;
	-- signal N3_19_34 : std_logic;
	HA28 : half_adder port map (N0_27_33,N0_28_33,N3_18_33,N3_19_34);
-- In matrix 2 adding FA to column 34 
	-- signal N3_0_34 : std_logic;
	-- signal N3_1_35 : std_logic;
	FA334 : full_adder port map (N0_0_34,N0_1_34,N0_2_34,N3_0_34,N3_1_35);
-- In matrix 2 adding FA to column 34 
	-- signal N3_2_34 : std_logic;
	-- signal N3_3_35 : std_logic;
	FA335 : full_adder port map (N0_3_34,N0_4_34,N0_5_34,N3_2_34,N3_3_35);
-- In matrix 2 adding FA to column 34 
	-- signal N3_4_34 : std_logic;
	-- signal N3_5_35 : std_logic;
	FA336 : full_adder port map (N0_6_34,N0_7_34,N0_8_34,N3_4_34,N3_5_35);
-- In matrix 2 adding FA to column 34 
	-- signal N3_6_34 : std_logic;
	-- signal N3_7_35 : std_logic;
	FA337 : full_adder port map (N0_9_34,N0_10_34,N0_11_34,N3_6_34,N3_7_35);
-- In matrix 2 adding FA to column 34 
	-- signal N3_8_34 : std_logic;
	-- signal N3_9_35 : std_logic;
	FA338 : full_adder port map (N0_12_34,N0_13_34,N0_14_34,N3_8_34,N3_9_35);
-- In matrix 2 adding FA to column 34 
	-- signal N3_10_34 : std_logic;
	-- signal N3_11_35 : std_logic;
	FA339 : full_adder port map (N0_15_34,N0_16_34,N0_17_34,N3_10_34,N3_11_35);
-- In matrix 2 adding FA to column 34 
	-- signal N3_12_34 : std_logic;
	-- signal N3_13_35 : std_logic;
	FA340 : full_adder port map (N0_18_34,N0_19_34,N0_20_34,N3_12_34,N3_13_35);
-- In matrix 2 adding FA to column 34 
	-- signal N3_14_34 : std_logic;
	-- signal N3_15_35 : std_logic;
	FA341 : full_adder port map (N0_21_34,N0_22_34,N0_23_34,N3_14_34,N3_15_35);
-- In matrix 2 adding FA to column 34 
	-- signal N3_16_34 : std_logic;
	-- signal N3_17_35 : std_logic;
	FA342 : full_adder port map (N0_24_34,N0_25_34,N0_26_34,N3_16_34,N3_17_35);
-- In matrix 2 adding FA to column 34 
	-- signal N3_18_34 : std_logic;
	-- signal N3_19_35 : std_logic;
	FA343 : full_adder port map (N0_27_34,N0_28_34,N0_29_34,N3_18_34,N3_19_35);
-- In matrix 2 adding HA to column 34 
	-- signal N3_20_34 : std_logic;
	-- signal N3_21_35 : std_logic;
	HA29 : half_adder port map (N0_30_34,N0_31_34,N3_20_34,N3_21_35);
-- In matrix 2 adding FA to column 35 
	-- signal N3_0_35 : std_logic;
	-- signal N3_1_36 : std_logic;
	FA344 : full_adder port map (N0_0_35,N0_1_35,N0_2_35,N3_0_35,N3_1_36);
-- In matrix 2 adding FA to column 35 
	-- signal N3_2_35 : std_logic;
	-- signal N3_3_36 : std_logic;
	FA345 : full_adder port map (N0_3_35,N0_4_35,N0_5_35,N3_2_35,N3_3_36);
-- In matrix 2 adding FA to column 35 
	-- signal N3_4_35 : std_logic;
	-- signal N3_5_36 : std_logic;
	FA346 : full_adder port map (N0_6_35,N0_7_35,N0_8_35,N3_4_35,N3_5_36);
-- In matrix 2 adding FA to column 35 
	-- signal N3_6_35 : std_logic;
	-- signal N3_7_36 : std_logic;
	FA347 : full_adder port map (N0_9_35,N0_10_35,N0_11_35,N3_6_35,N3_7_36);
-- In matrix 2 adding FA to column 35 
	-- signal N3_8_35 : std_logic;
	-- signal N3_9_36 : std_logic;
	FA348 : full_adder port map (N0_12_35,N0_13_35,N0_14_35,N3_8_35,N3_9_36);
-- In matrix 2 adding FA to column 35 
	-- signal N3_10_35 : std_logic;
	-- signal N3_11_36 : std_logic;
	FA349 : full_adder port map (N0_15_35,N0_16_35,N0_17_35,N3_10_35,N3_11_36);
-- In matrix 2 adding FA to column 35 
	-- signal N3_12_35 : std_logic;
	-- signal N3_13_36 : std_logic;
	FA350 : full_adder port map (N0_18_35,N0_19_35,N0_20_35,N3_12_35,N3_13_36);
-- In matrix 2 adding FA to column 35 
	-- signal N3_14_35 : std_logic;
	-- signal N3_15_36 : std_logic;
	FA351 : full_adder port map (N0_21_35,N0_22_35,N0_23_35,N3_14_35,N3_15_36);
-- In matrix 2 adding FA to column 35 
	-- signal N3_16_35 : std_logic;
	-- signal N3_17_36 : std_logic;
	FA352 : full_adder port map (N0_24_35,N0_25_35,N0_26_35,N3_16_35,N3_17_36);
-- In matrix 2 adding FA to column 35 
	-- signal N3_18_35 : std_logic;
	-- signal N3_19_36 : std_logic;
	FA353 : full_adder port map (N0_27_35,N0_28_35,N0_29_35,N3_18_35,N3_19_36);
-- In matrix 2 adding FA to column 35 
	-- signal N3_20_35 : std_logic;
	-- signal N3_21_36 : std_logic;
	FA354 : full_adder port map (N0_30_35,N0_31_35,N0_32_35,N3_20_35,N3_21_36);
-- In matrix 2 adding HA to column 35 
	-- signal N3_22_35 : std_logic;
	-- signal N3_23_36 : std_logic;
	HA30 : half_adder port map (N0_33_35,N0_34_35,N3_22_35,N3_23_36);
-- In matrix 2 adding FA to column 36 
	-- signal N3_0_36 : std_logic;
	-- signal N3_1_37 : std_logic;
	FA355 : full_adder port map (N0_2_36,N0_3_36,N0_4_36,N3_0_36,N3_1_37);
-- In matrix 2 adding FA to column 36 
	-- signal N3_2_36 : std_logic;
	-- signal N3_3_37 : std_logic;
	FA356 : full_adder port map (N0_5_36,N0_6_36,N0_7_36,N3_2_36,N3_3_37);
-- In matrix 2 adding FA to column 36 
	-- signal N3_4_36 : std_logic;
	-- signal N3_5_37 : std_logic;
	FA357 : full_adder port map (N0_8_36,N0_9_36,N0_10_36,N3_4_36,N3_5_37);
-- In matrix 2 adding FA to column 36 
	-- signal N3_6_36 : std_logic;
	-- signal N3_7_37 : std_logic;
	FA358 : full_adder port map (N0_11_36,N0_12_36,N0_13_36,N3_6_36,N3_7_37);
-- In matrix 2 adding FA to column 36 
	-- signal N3_8_36 : std_logic;
	-- signal N3_9_37 : std_logic;
	FA359 : full_adder port map (N0_14_36,N0_15_36,N0_16_36,N3_8_36,N3_9_37);
-- In matrix 2 adding FA to column 36 
	-- signal N3_10_36 : std_logic;
	-- signal N3_11_37 : std_logic;
	FA360 : full_adder port map (N0_17_36,N0_18_36,N0_19_36,N3_10_36,N3_11_37);
-- In matrix 2 adding FA to column 36 
	-- signal N3_12_36 : std_logic;
	-- signal N3_13_37 : std_logic;
	FA361 : full_adder port map (N0_20_36,N0_21_36,N0_22_36,N3_12_36,N3_13_37);
-- In matrix 2 adding FA to column 36 
	-- signal N3_14_36 : std_logic;
	-- signal N3_15_37 : std_logic;
	FA362 : full_adder port map (N0_23_36,N0_24_36,N0_25_36,N3_14_36,N3_15_37);
-- In matrix 2 adding FA to column 36 
	-- signal N3_16_36 : std_logic;
	-- signal N3_17_37 : std_logic;
	FA363 : full_adder port map (N0_26_36,N0_27_36,N0_28_36,N3_16_36,N3_17_37);
-- In matrix 2 adding FA to column 36 
	-- signal N3_18_36 : std_logic;
	-- signal N3_19_37 : std_logic;
	FA364 : full_adder port map (N0_29_36,N0_30_36,N0_31_36,N3_18_36,N3_19_37);
-- In matrix 2 adding FA to column 36 
	-- signal N3_20_36 : std_logic;
	-- signal N3_21_37 : std_logic;
	FA365 : full_adder port map (N0_32_36,N0_33_36,N0_34_36,N3_20_36,N3_21_37);
-- In matrix 2 adding FA to column 36 
	-- signal N3_22_36 : std_logic;
	-- signal N3_23_37 : std_logic;
	FA366 : full_adder port map (N0_35_36,N0_36_36,N2_0_36,N3_22_36,N3_23_37);
-- In matrix 2 adding FA to column 37 
	-- signal N3_0_37 : std_logic;
	-- signal N3_1_38 : std_logic;
	FA367 : full_adder port map (N0_5_37,N0_6_37,N0_7_37,N3_0_37,N3_1_38);
-- In matrix 2 adding FA to column 37 
	-- signal N3_2_37 : std_logic;
	-- signal N3_3_38 : std_logic;
	FA368 : full_adder port map (N0_8_37,N0_9_37,N0_10_37,N3_2_37,N3_3_38);
-- In matrix 2 adding FA to column 37 
	-- signal N3_4_37 : std_logic;
	-- signal N3_5_38 : std_logic;
	FA369 : full_adder port map (N0_11_37,N0_12_37,N0_13_37,N3_4_37,N3_5_38);
-- In matrix 2 adding FA to column 37 
	-- signal N3_6_37 : std_logic;
	-- signal N3_7_38 : std_logic;
	FA370 : full_adder port map (N0_14_37,N0_15_37,N0_16_37,N3_6_37,N3_7_38);
-- In matrix 2 adding FA to column 37 
	-- signal N3_8_37 : std_logic;
	-- signal N3_9_38 : std_logic;
	FA371 : full_adder port map (N0_17_37,N0_18_37,N0_19_37,N3_8_37,N3_9_38);
-- In matrix 2 adding FA to column 37 
	-- signal N3_10_37 : std_logic;
	-- signal N3_11_38 : std_logic;
	FA372 : full_adder port map (N0_20_37,N0_21_37,N0_22_37,N3_10_37,N3_11_38);
-- In matrix 2 adding FA to column 37 
	-- signal N3_12_37 : std_logic;
	-- signal N3_13_38 : std_logic;
	FA373 : full_adder port map (N0_23_37,N0_24_37,N0_25_37,N3_12_37,N3_13_38);
-- In matrix 2 adding FA to column 37 
	-- signal N3_14_37 : std_logic;
	-- signal N3_15_38 : std_logic;
	FA374 : full_adder port map (N0_26_37,N0_27_37,N0_28_37,N3_14_37,N3_15_38);
-- In matrix 2 adding FA to column 37 
	-- signal N3_16_37 : std_logic;
	-- signal N3_17_38 : std_logic;
	FA375 : full_adder port map (N0_29_37,N0_30_37,N0_31_37,N3_16_37,N3_17_38);
-- In matrix 2 adding FA to column 37 
	-- signal N3_18_37 : std_logic;
	-- signal N3_19_38 : std_logic;
	FA376 : full_adder port map (N0_32_37,N0_33_37,N0_34_37,N3_18_37,N3_19_38);
-- In matrix 2 adding FA to column 37 
	-- signal N3_20_37 : std_logic;
	-- signal N3_21_38 : std_logic;
	FA377 : full_adder port map (N0_35_37,N0_36_37,N0_37_37,N3_20_37,N3_21_38);
-- In matrix 2 adding FA to column 37 
	-- signal N3_22_37 : std_logic;
	-- signal N3_23_38 : std_logic;
	FA378 : full_adder port map (N2_0_37,N2_1_37,N2_2_37,N3_22_37,N3_23_38);
-- In matrix 2 adding FA to column 38 
	-- signal N3_0_38 : std_logic;
	-- signal N3_1_39 : std_logic;
	FA379 : full_adder port map (N0_8_38,N0_9_38,N0_10_38,N3_0_38,N3_1_39);
-- In matrix 2 adding FA to column 38 
	-- signal N3_2_38 : std_logic;
	-- signal N3_3_39 : std_logic;
	FA380 : full_adder port map (N0_11_38,N0_12_38,N0_13_38,N3_2_38,N3_3_39);
-- In matrix 2 adding FA to column 38 
	-- signal N3_4_38 : std_logic;
	-- signal N3_5_39 : std_logic;
	FA381 : full_adder port map (N0_14_38,N0_15_38,N0_16_38,N3_4_38,N3_5_39);
-- In matrix 2 adding FA to column 38 
	-- signal N3_6_38 : std_logic;
	-- signal N3_7_39 : std_logic;
	FA382 : full_adder port map (N0_17_38,N0_18_38,N0_19_38,N3_6_38,N3_7_39);
-- In matrix 2 adding FA to column 38 
	-- signal N3_8_38 : std_logic;
	-- signal N3_9_39 : std_logic;
	FA383 : full_adder port map (N0_20_38,N0_21_38,N0_22_38,N3_8_38,N3_9_39);
-- In matrix 2 adding FA to column 38 
	-- signal N3_10_38 : std_logic;
	-- signal N3_11_39 : std_logic;
	FA384 : full_adder port map (N0_23_38,N0_24_38,N0_25_38,N3_10_38,N3_11_39);
-- In matrix 2 adding FA to column 38 
	-- signal N3_12_38 : std_logic;
	-- signal N3_13_39 : std_logic;
	FA385 : full_adder port map (N0_26_38,N0_27_38,N0_28_38,N3_12_38,N3_13_39);
-- In matrix 2 adding FA to column 38 
	-- signal N3_14_38 : std_logic;
	-- signal N3_15_39 : std_logic;
	FA386 : full_adder port map (N0_29_38,N0_30_38,N0_31_38,N3_14_38,N3_15_39);
-- In matrix 2 adding FA to column 38 
	-- signal N3_16_38 : std_logic;
	-- signal N3_17_39 : std_logic;
	FA387 : full_adder port map (N0_32_38,N0_33_38,N0_34_38,N3_16_38,N3_17_39);
-- In matrix 2 adding FA to column 38 
	-- signal N3_18_38 : std_logic;
	-- signal N3_19_39 : std_logic;
	FA388 : full_adder port map (N0_35_38,N0_36_38,N0_37_38,N3_18_38,N3_19_39);
-- In matrix 2 adding FA to column 38 
	-- signal N3_20_38 : std_logic;
	-- signal N3_21_39 : std_logic;
	FA389 : full_adder port map (N0_38_38,N2_0_38,N2_1_38,N3_20_38,N3_21_39);
-- In matrix 2 adding FA to column 38 
	-- signal N3_22_38 : std_logic;
	-- signal N3_23_39 : std_logic;
	FA390 : full_adder port map (N2_2_38,N2_3_38,N2_4_38,N3_22_38,N3_23_39);
-- In matrix 2 adding FA to column 39 
	-- signal N3_0_39 : std_logic;
	-- signal N3_1_40 : std_logic;
	FA391 : full_adder port map (N0_11_39,N0_12_39,N0_13_39,N3_0_39,N3_1_40);
-- In matrix 2 adding FA to column 39 
	-- signal N3_2_39 : std_logic;
	-- signal N3_3_40 : std_logic;
	FA392 : full_adder port map (N0_14_39,N0_15_39,N0_16_39,N3_2_39,N3_3_40);
-- In matrix 2 adding FA to column 39 
	-- signal N3_4_39 : std_logic;
	-- signal N3_5_40 : std_logic;
	FA393 : full_adder port map (N0_17_39,N0_18_39,N0_19_39,N3_4_39,N3_5_40);
-- In matrix 2 adding FA to column 39 
	-- signal N3_6_39 : std_logic;
	-- signal N3_7_40 : std_logic;
	FA394 : full_adder port map (N0_20_39,N0_21_39,N0_22_39,N3_6_39,N3_7_40);
-- In matrix 2 adding FA to column 39 
	-- signal N3_8_39 : std_logic;
	-- signal N3_9_40 : std_logic;
	FA395 : full_adder port map (N0_23_39,N0_24_39,N0_25_39,N3_8_39,N3_9_40);
-- In matrix 2 adding FA to column 39 
	-- signal N3_10_39 : std_logic;
	-- signal N3_11_40 : std_logic;
	FA396 : full_adder port map (N0_26_39,N0_27_39,N0_28_39,N3_10_39,N3_11_40);
-- In matrix 2 adding FA to column 39 
	-- signal N3_12_39 : std_logic;
	-- signal N3_13_40 : std_logic;
	FA397 : full_adder port map (N0_29_39,N0_30_39,N0_31_39,N3_12_39,N3_13_40);
-- In matrix 2 adding FA to column 39 
	-- signal N3_14_39 : std_logic;
	-- signal N3_15_40 : std_logic;
	FA398 : full_adder port map (N0_32_39,N0_33_39,N0_34_39,N3_14_39,N3_15_40);
-- In matrix 2 adding FA to column 39 
	-- signal N3_16_39 : std_logic;
	-- signal N3_17_40 : std_logic;
	FA399 : full_adder port map (N0_35_39,N0_36_39,N0_37_39,N3_16_39,N3_17_40);
-- In matrix 2 adding FA to column 39 
	-- signal N3_18_39 : std_logic;
	-- signal N3_19_40 : std_logic;
	FA400 : full_adder port map (N0_38_39,N0_39_39,N2_0_39,N3_18_39,N3_19_40);
-- In matrix 2 adding FA to column 39 
	-- signal N3_20_39 : std_logic;
	-- signal N3_21_40 : std_logic;
	FA401 : full_adder port map (N2_1_39,N2_2_39,N2_3_39,N3_20_39,N3_21_40);
-- In matrix 2 adding FA to column 39 
	-- signal N3_22_39 : std_logic;
	-- signal N3_23_40 : std_logic;
	FA402 : full_adder port map (N2_4_39,N2_5_39,N2_6_39,N3_22_39,N3_23_40);
-- In matrix 2 adding FA to column 40 
	-- signal N3_0_40 : std_logic;
	-- signal N3_1_41 : std_logic;
	FA403 : full_adder port map (N0_14_40,N0_15_40,N0_16_40,N3_0_40,N3_1_41);
-- In matrix 2 adding FA to column 40 
	-- signal N3_2_40 : std_logic;
	-- signal N3_3_41 : std_logic;
	FA404 : full_adder port map (N0_17_40,N0_18_40,N0_19_40,N3_2_40,N3_3_41);
-- In matrix 2 adding FA to column 40 
	-- signal N3_4_40 : std_logic;
	-- signal N3_5_41 : std_logic;
	FA405 : full_adder port map (N0_20_40,N0_21_40,N0_22_40,N3_4_40,N3_5_41);
-- In matrix 2 adding FA to column 40 
	-- signal N3_6_40 : std_logic;
	-- signal N3_7_41 : std_logic;
	FA406 : full_adder port map (N0_23_40,N0_24_40,N0_25_40,N3_6_40,N3_7_41);
-- In matrix 2 adding FA to column 40 
	-- signal N3_8_40 : std_logic;
	-- signal N3_9_41 : std_logic;
	FA407 : full_adder port map (N0_26_40,N0_27_40,N0_28_40,N3_8_40,N3_9_41);
-- In matrix 2 adding FA to column 40 
	-- signal N3_10_40 : std_logic;
	-- signal N3_11_41 : std_logic;
	FA408 : full_adder port map (N0_29_40,N0_30_40,N0_31_40,N3_10_40,N3_11_41);
-- In matrix 2 adding FA to column 40 
	-- signal N3_12_40 : std_logic;
	-- signal N3_13_41 : std_logic;
	FA409 : full_adder port map (N0_32_40,N0_33_40,N0_34_40,N3_12_40,N3_13_41);
-- In matrix 2 adding FA to column 40 
	-- signal N3_14_40 : std_logic;
	-- signal N3_15_41 : std_logic;
	FA410 : full_adder port map (N0_35_40,N0_36_40,N0_37_40,N3_14_40,N3_15_41);
-- In matrix 2 adding FA to column 40 
	-- signal N3_16_40 : std_logic;
	-- signal N3_17_41 : std_logic;
	FA411 : full_adder port map (N0_38_40,N0_39_40,N0_40_40,N3_16_40,N3_17_41);
-- In matrix 2 adding FA to column 40 
	-- signal N3_18_40 : std_logic;
	-- signal N3_19_41 : std_logic;
	FA412 : full_adder port map (N2_0_40,N2_1_40,N2_2_40,N3_18_40,N3_19_41);
-- In matrix 2 adding FA to column 40 
	-- signal N3_20_40 : std_logic;
	-- signal N3_21_41 : std_logic;
	FA413 : full_adder port map (N2_3_40,N2_4_40,N2_5_40,N3_20_40,N3_21_41);
-- In matrix 2 adding FA to column 40 
	-- signal N3_22_40 : std_logic;
	-- signal N3_23_41 : std_logic;
	FA414 : full_adder port map (N2_6_40,N2_7_40,N2_8_40,N3_22_40,N3_23_41);
-- In matrix 2 adding FA to column 41 
	-- signal N3_0_41 : std_logic;
	-- signal N3_1_42 : std_logic;
	FA415 : full_adder port map (N0_17_41,N0_18_41,N0_19_41,N3_0_41,N3_1_42);
-- In matrix 2 adding FA to column 41 
	-- signal N3_2_41 : std_logic;
	-- signal N3_3_42 : std_logic;
	FA416 : full_adder port map (N0_20_41,N0_21_41,N0_22_41,N3_2_41,N3_3_42);
-- In matrix 2 adding FA to column 41 
	-- signal N3_4_41 : std_logic;
	-- signal N3_5_42 : std_logic;
	FA417 : full_adder port map (N0_23_41,N0_24_41,N0_25_41,N3_4_41,N3_5_42);
-- In matrix 2 adding FA to column 41 
	-- signal N3_6_41 : std_logic;
	-- signal N3_7_42 : std_logic;
	FA418 : full_adder port map (N0_26_41,N0_27_41,N0_28_41,N3_6_41,N3_7_42);
-- In matrix 2 adding FA to column 41 
	-- signal N3_8_41 : std_logic;
	-- signal N3_9_42 : std_logic;
	FA419 : full_adder port map (N0_29_41,N0_30_41,N0_31_41,N3_8_41,N3_9_42);
-- In matrix 2 adding FA to column 41 
	-- signal N3_10_41 : std_logic;
	-- signal N3_11_42 : std_logic;
	FA420 : full_adder port map (N0_32_41,N0_33_41,N0_34_41,N3_10_41,N3_11_42);
-- In matrix 2 adding FA to column 41 
	-- signal N3_12_41 : std_logic;
	-- signal N3_13_42 : std_logic;
	FA421 : full_adder port map (N0_35_41,N0_36_41,N0_37_41,N3_12_41,N3_13_42);
-- In matrix 2 adding FA to column 41 
	-- signal N3_14_41 : std_logic;
	-- signal N3_15_42 : std_logic;
	FA422 : full_adder port map (N0_38_41,N0_39_41,N0_40_41,N3_14_41,N3_15_42);
-- In matrix 2 adding FA to column 41 
	-- signal N3_16_41 : std_logic;
	-- signal N3_17_42 : std_logic;
	FA423 : full_adder port map (N0_41_41,N2_0_41,N2_1_41,N3_16_41,N3_17_42);
-- In matrix 2 adding FA to column 41 
	-- signal N3_18_41 : std_logic;
	-- signal N3_19_42 : std_logic;
	FA424 : full_adder port map (N2_2_41,N2_3_41,N2_4_41,N3_18_41,N3_19_42);
-- In matrix 2 adding FA to column 41 
	-- signal N3_20_41 : std_logic;
	-- signal N3_21_42 : std_logic;
	FA425 : full_adder port map (N2_5_41,N2_6_41,N2_7_41,N3_20_41,N3_21_42);
-- In matrix 2 adding FA to column 41 
	-- signal N3_22_41 : std_logic;
	-- signal N3_23_42 : std_logic;
	FA426 : full_adder port map (N2_8_41,N2_9_41,N2_10_41,N3_22_41,N3_23_42);
-- In matrix 2 adding FA to column 42 
	-- signal N3_0_42 : std_logic;
	-- signal N3_1_43 : std_logic;
	FA427 : full_adder port map (N0_20_42,N0_21_42,N0_22_42,N3_0_42,N3_1_43);
-- In matrix 2 adding FA to column 42 
	-- signal N3_2_42 : std_logic;
	-- signal N3_3_43 : std_logic;
	FA428 : full_adder port map (N0_23_42,N0_24_42,N0_25_42,N3_2_42,N3_3_43);
-- In matrix 2 adding FA to column 42 
	-- signal N3_4_42 : std_logic;
	-- signal N3_5_43 : std_logic;
	FA429 : full_adder port map (N0_26_42,N0_27_42,N0_28_42,N3_4_42,N3_5_43);
-- In matrix 2 adding FA to column 42 
	-- signal N3_6_42 : std_logic;
	-- signal N3_7_43 : std_logic;
	FA430 : full_adder port map (N0_29_42,N0_30_42,N0_31_42,N3_6_42,N3_7_43);
-- In matrix 2 adding FA to column 42 
	-- signal N3_8_42 : std_logic;
	-- signal N3_9_43 : std_logic;
	FA431 : full_adder port map (N0_32_42,N0_33_42,N0_34_42,N3_8_42,N3_9_43);
-- In matrix 2 adding FA to column 42 
	-- signal N3_10_42 : std_logic;
	-- signal N3_11_43 : std_logic;
	FA432 : full_adder port map (N0_35_42,N0_36_42,N0_37_42,N3_10_42,N3_11_43);
-- In matrix 2 adding FA to column 42 
	-- signal N3_12_42 : std_logic;
	-- signal N3_13_43 : std_logic;
	FA433 : full_adder port map (N0_38_42,N0_39_42,N0_40_42,N3_12_42,N3_13_43);
-- In matrix 2 adding FA to column 42 
	-- signal N3_14_42 : std_logic;
	-- signal N3_15_43 : std_logic;
	FA434 : full_adder port map (N0_41_42,N0_42_42,N2_0_42,N3_14_42,N3_15_43);
-- In matrix 2 adding FA to column 42 
	-- signal N3_16_42 : std_logic;
	-- signal N3_17_43 : std_logic;
	FA435 : full_adder port map (N2_1_42,N2_2_42,N2_3_42,N3_16_42,N3_17_43);
-- In matrix 2 adding FA to column 42 
	-- signal N3_18_42 : std_logic;
	-- signal N3_19_43 : std_logic;
	FA436 : full_adder port map (N2_4_42,N2_5_42,N2_6_42,N3_18_42,N3_19_43);
-- In matrix 2 adding FA to column 42 
	-- signal N3_20_42 : std_logic;
	-- signal N3_21_43 : std_logic;
	FA437 : full_adder port map (N2_7_42,N2_8_42,N2_9_42,N3_20_42,N3_21_43);
-- In matrix 2 adding FA to column 42 
	-- signal N3_22_42 : std_logic;
	-- signal N3_23_43 : std_logic;
	FA438 : full_adder port map (N2_10_42,N2_11_42,N2_12_42,N3_22_42,N3_23_43);
-- In matrix 2 adding FA to column 43 
	-- signal N3_0_43 : std_logic;
	-- signal N3_1_44 : std_logic;
	FA439 : full_adder port map (N0_23_43,N0_24_43,N0_25_43,N3_0_43,N3_1_44);
-- In matrix 2 adding FA to column 43 
	-- signal N3_2_43 : std_logic;
	-- signal N3_3_44 : std_logic;
	FA440 : full_adder port map (N0_26_43,N0_27_43,N0_28_43,N3_2_43,N3_3_44);
-- In matrix 2 adding FA to column 43 
	-- signal N3_4_43 : std_logic;
	-- signal N3_5_44 : std_logic;
	FA441 : full_adder port map (N0_29_43,N0_30_43,N0_31_43,N3_4_43,N3_5_44);
-- In matrix 2 adding FA to column 43 
	-- signal N3_6_43 : std_logic;
	-- signal N3_7_44 : std_logic;
	FA442 : full_adder port map (N0_32_43,N0_33_43,N0_34_43,N3_6_43,N3_7_44);
-- In matrix 2 adding FA to column 43 
	-- signal N3_8_43 : std_logic;
	-- signal N3_9_44 : std_logic;
	FA443 : full_adder port map (N0_35_43,N0_36_43,N0_37_43,N3_8_43,N3_9_44);
-- In matrix 2 adding FA to column 43 
	-- signal N3_10_43 : std_logic;
	-- signal N3_11_44 : std_logic;
	FA444 : full_adder port map (N0_38_43,N0_39_43,N0_40_43,N3_10_43,N3_11_44);
-- In matrix 2 adding FA to column 43 
	-- signal N3_12_43 : std_logic;
	-- signal N3_13_44 : std_logic;
	FA445 : full_adder port map (N0_41_43,N0_42_43,N0_43_43,N3_12_43,N3_13_44);
-- In matrix 2 adding FA to column 43 
	-- signal N3_14_43 : std_logic;
	-- signal N3_15_44 : std_logic;
	FA446 : full_adder port map (N2_0_43,N2_1_43,N2_2_43,N3_14_43,N3_15_44);
-- In matrix 2 adding FA to column 43 
	-- signal N3_16_43 : std_logic;
	-- signal N3_17_44 : std_logic;
	FA447 : full_adder port map (N2_3_43,N2_4_43,N2_5_43,N3_16_43,N3_17_44);
-- In matrix 2 adding FA to column 43 
	-- signal N3_18_43 : std_logic;
	-- signal N3_19_44 : std_logic;
	FA448 : full_adder port map (N2_6_43,N2_7_43,N2_8_43,N3_18_43,N3_19_44);
-- In matrix 2 adding FA to column 43 
	-- signal N3_20_43 : std_logic;
	-- signal N3_21_44 : std_logic;
	FA449 : full_adder port map (N2_9_43,N2_10_43,N2_11_43,N3_20_43,N3_21_44);
-- In matrix 2 adding FA to column 43 
	-- signal N3_22_43 : std_logic;
	-- signal N3_23_44 : std_logic;
	FA450 : full_adder port map (N2_12_43,N2_13_43,N2_14_43,N3_22_43,N3_23_44);
-- In matrix 2 adding FA to column 44 
	-- signal N3_0_44 : std_logic;
	-- signal N3_1_45 : std_logic;
	FA451 : full_adder port map (N0_26_44,N0_27_44,N0_28_44,N3_0_44,N3_1_45);
-- In matrix 2 adding FA to column 44 
	-- signal N3_2_44 : std_logic;
	-- signal N3_3_45 : std_logic;
	FA452 : full_adder port map (N0_29_44,N0_30_44,N0_31_44,N3_2_44,N3_3_45);
-- In matrix 2 adding FA to column 44 
	-- signal N3_4_44 : std_logic;
	-- signal N3_5_45 : std_logic;
	FA453 : full_adder port map (N0_32_44,N0_33_44,N0_34_44,N3_4_44,N3_5_45);
-- In matrix 2 adding FA to column 44 
	-- signal N3_6_44 : std_logic;
	-- signal N3_7_45 : std_logic;
	FA454 : full_adder port map (N0_35_44,N0_36_44,N0_37_44,N3_6_44,N3_7_45);
-- In matrix 2 adding FA to column 44 
	-- signal N3_8_44 : std_logic;
	-- signal N3_9_45 : std_logic;
	FA455 : full_adder port map (N0_38_44,N0_39_44,N0_40_44,N3_8_44,N3_9_45);
-- In matrix 2 adding FA to column 44 
	-- signal N3_10_44 : std_logic;
	-- signal N3_11_45 : std_logic;
	FA456 : full_adder port map (N0_41_44,N0_42_44,N0_43_44,N3_10_44,N3_11_45);
-- In matrix 2 adding FA to column 44 
	-- signal N3_12_44 : std_logic;
	-- signal N3_13_45 : std_logic;
	FA457 : full_adder port map (N0_44_44,N2_0_44,N2_1_44,N3_12_44,N3_13_45);
-- In matrix 2 adding FA to column 44 
	-- signal N3_14_44 : std_logic;
	-- signal N3_15_45 : std_logic;
	FA458 : full_adder port map (N2_2_44,N2_3_44,N2_4_44,N3_14_44,N3_15_45);
-- In matrix 2 adding FA to column 44 
	-- signal N3_16_44 : std_logic;
	-- signal N3_17_45 : std_logic;
	FA459 : full_adder port map (N2_5_44,N2_6_44,N2_7_44,N3_16_44,N3_17_45);
-- In matrix 2 adding FA to column 44 
	-- signal N3_18_44 : std_logic;
	-- signal N3_19_45 : std_logic;
	FA460 : full_adder port map (N2_8_44,N2_9_44,N2_10_44,N3_18_44,N3_19_45);
-- In matrix 2 adding FA to column 44 
	-- signal N3_20_44 : std_logic;
	-- signal N3_21_45 : std_logic;
	FA461 : full_adder port map (N2_11_44,N2_12_44,N2_13_44,N3_20_44,N3_21_45);
-- In matrix 2 adding FA to column 44 
	-- signal N3_22_44 : std_logic;
	-- signal N3_23_45 : std_logic;
	FA462 : full_adder port map (N2_14_44,N2_15_44,N2_16_44,N3_22_44,N3_23_45);
-- In matrix 2 adding FA to column 45 
	-- signal N3_0_45 : std_logic;
	-- signal N3_1_46 : std_logic;
	FA463 : full_adder port map (N0_29_45,N0_30_45,N0_31_45,N3_0_45,N3_1_46);
-- In matrix 2 adding FA to column 45 
	-- signal N3_2_45 : std_logic;
	-- signal N3_3_46 : std_logic;
	FA464 : full_adder port map (N0_32_45,N0_33_45,N0_34_45,N3_2_45,N3_3_46);
-- In matrix 2 adding FA to column 45 
	-- signal N3_4_45 : std_logic;
	-- signal N3_5_46 : std_logic;
	FA465 : full_adder port map (N0_35_45,N0_36_45,N0_37_45,N3_4_45,N3_5_46);
-- In matrix 2 adding FA to column 45 
	-- signal N3_6_45 : std_logic;
	-- signal N3_7_46 : std_logic;
	FA466 : full_adder port map (N0_38_45,N0_39_45,N0_40_45,N3_6_45,N3_7_46);
-- In matrix 2 adding FA to column 45 
	-- signal N3_8_45 : std_logic;
	-- signal N3_9_46 : std_logic;
	FA467 : full_adder port map (N0_41_45,N0_42_45,N0_43_45,N3_8_45,N3_9_46);
-- In matrix 2 adding FA to column 45 
	-- signal N3_10_45 : std_logic;
	-- signal N3_11_46 : std_logic;
	FA468 : full_adder port map (N0_44_45,N0_45_45,N2_0_45,N3_10_45,N3_11_46);
-- In matrix 2 adding FA to column 45 
	-- signal N3_12_45 : std_logic;
	-- signal N3_13_46 : std_logic;
	FA469 : full_adder port map (N2_1_45,N2_2_45,N2_3_45,N3_12_45,N3_13_46);
-- In matrix 2 adding FA to column 45 
	-- signal N3_14_45 : std_logic;
	-- signal N3_15_46 : std_logic;
	FA470 : full_adder port map (N2_4_45,N2_5_45,N2_6_45,N3_14_45,N3_15_46);
-- In matrix 2 adding FA to column 45 
	-- signal N3_16_45 : std_logic;
	-- signal N3_17_46 : std_logic;
	FA471 : full_adder port map (N2_7_45,N2_8_45,N2_9_45,N3_16_45,N3_17_46);
-- In matrix 2 adding FA to column 45 
	-- signal N3_18_45 : std_logic;
	-- signal N3_19_46 : std_logic;
	FA472 : full_adder port map (N2_10_45,N2_11_45,N2_12_45,N3_18_45,N3_19_46);
-- In matrix 2 adding FA to column 45 
	-- signal N3_20_45 : std_logic;
	-- signal N3_21_46 : std_logic;
	FA473 : full_adder port map (N2_13_45,N2_14_45,N2_15_45,N3_20_45,N3_21_46);
-- In matrix 2 adding FA to column 45 
	-- signal N3_22_45 : std_logic;
	-- signal N3_23_46 : std_logic;
	FA474 : full_adder port map (N2_16_45,N2_17_45,N2_18_45,N3_22_45,N3_23_46);
-- In matrix 2 adding FA to column 46 
	-- signal N3_0_46 : std_logic;
	-- signal N3_1_47 : std_logic;
	FA475 : full_adder port map (N0_32_46,N0_33_46,N0_34_46,N3_0_46,N3_1_47);
-- In matrix 2 adding FA to column 46 
	-- signal N3_2_46 : std_logic;
	-- signal N3_3_47 : std_logic;
	FA476 : full_adder port map (N0_35_46,N0_36_46,N0_37_46,N3_2_46,N3_3_47);
-- In matrix 2 adding FA to column 46 
	-- signal N3_4_46 : std_logic;
	-- signal N3_5_47 : std_logic;
	FA477 : full_adder port map (N0_38_46,N0_39_46,N0_40_46,N3_4_46,N3_5_47);
-- In matrix 2 adding FA to column 46 
	-- signal N3_6_46 : std_logic;
	-- signal N3_7_47 : std_logic;
	FA478 : full_adder port map (N0_41_46,N0_42_46,N0_43_46,N3_6_46,N3_7_47);
-- In matrix 2 adding FA to column 46 
	-- signal N3_8_46 : std_logic;
	-- signal N3_9_47 : std_logic;
	FA479 : full_adder port map (N0_44_46,N0_45_46,N0_46_46,N3_8_46,N3_9_47);
-- In matrix 2 adding FA to column 46 
	-- signal N3_10_46 : std_logic;
	-- signal N3_11_47 : std_logic;
	FA480 : full_adder port map (N2_0_46,N2_1_46,N2_2_46,N3_10_46,N3_11_47);
-- In matrix 2 adding FA to column 46 
	-- signal N3_12_46 : std_logic;
	-- signal N3_13_47 : std_logic;
	FA481 : full_adder port map (N2_3_46,N2_4_46,N2_5_46,N3_12_46,N3_13_47);
-- In matrix 2 adding FA to column 46 
	-- signal N3_14_46 : std_logic;
	-- signal N3_15_47 : std_logic;
	FA482 : full_adder port map (N2_6_46,N2_7_46,N2_8_46,N3_14_46,N3_15_47);
-- In matrix 2 adding FA to column 46 
	-- signal N3_16_46 : std_logic;
	-- signal N3_17_47 : std_logic;
	FA483 : full_adder port map (N2_9_46,N2_10_46,N2_11_46,N3_16_46,N3_17_47);
-- In matrix 2 adding FA to column 46 
	-- signal N3_18_46 : std_logic;
	-- signal N3_19_47 : std_logic;
	FA484 : full_adder port map (N2_12_46,N2_13_46,N2_14_46,N3_18_46,N3_19_47);
-- In matrix 2 adding FA to column 46 
	-- signal N3_20_46 : std_logic;
	-- signal N3_21_47 : std_logic;
	FA485 : full_adder port map (N2_15_46,N2_16_46,N2_17_46,N3_20_46,N3_21_47);
-- In matrix 2 adding FA to column 46 
	-- signal N3_22_46 : std_logic;
	-- signal N3_23_47 : std_logic;
	FA486 : full_adder port map (N2_18_46,N2_19_46,N2_20_46,N3_22_46,N3_23_47);
-- In matrix 2 adding FA to column 47 
	-- signal N3_0_47 : std_logic;
	-- signal N3_1_48 : std_logic;
	FA487 : full_adder port map (N0_35_47,N0_36_47,N0_37_47,N3_0_47,N3_1_48);
-- In matrix 2 adding FA to column 47 
	-- signal N3_2_47 : std_logic;
	-- signal N3_3_48 : std_logic;
	FA488 : full_adder port map (N0_38_47,N0_39_47,N0_40_47,N3_2_47,N3_3_48);
-- In matrix 2 adding FA to column 47 
	-- signal N3_4_47 : std_logic;
	-- signal N3_5_48 : std_logic;
	FA489 : full_adder port map (N0_41_47,N0_42_47,N0_43_47,N3_4_47,N3_5_48);
-- In matrix 2 adding FA to column 47 
	-- signal N3_6_47 : std_logic;
	-- signal N3_7_48 : std_logic;
	FA490 : full_adder port map (N0_44_47,N0_45_47,N0_46_47,N3_6_47,N3_7_48);
-- In matrix 2 adding FA to column 47 
	-- signal N3_8_47 : std_logic;
	-- signal N3_9_48 : std_logic;
	FA491 : full_adder port map (N0_47_47,N2_0_47,N2_1_47,N3_8_47,N3_9_48);
-- In matrix 2 adding FA to column 47 
	-- signal N3_10_47 : std_logic;
	-- signal N3_11_48 : std_logic;
	FA492 : full_adder port map (N2_2_47,N2_3_47,N2_4_47,N3_10_47,N3_11_48);
-- In matrix 2 adding FA to column 47 
	-- signal N3_12_47 : std_logic;
	-- signal N3_13_48 : std_logic;
	FA493 : full_adder port map (N2_5_47,N2_6_47,N2_7_47,N3_12_47,N3_13_48);
-- In matrix 2 adding FA to column 47 
	-- signal N3_14_47 : std_logic;
	-- signal N3_15_48 : std_logic;
	FA494 : full_adder port map (N2_8_47,N2_9_47,N2_10_47,N3_14_47,N3_15_48);
-- In matrix 2 adding FA to column 47 
	-- signal N3_16_47 : std_logic;
	-- signal N3_17_48 : std_logic;
	FA495 : full_adder port map (N2_11_47,N2_12_47,N2_13_47,N3_16_47,N3_17_48);
-- In matrix 2 adding FA to column 47 
	-- signal N3_18_47 : std_logic;
	-- signal N3_19_48 : std_logic;
	FA496 : full_adder port map (N2_14_47,N2_15_47,N2_16_47,N3_18_47,N3_19_48);
-- In matrix 2 adding FA to column 47 
	-- signal N3_20_47 : std_logic;
	-- signal N3_21_48 : std_logic;
	FA497 : full_adder port map (N2_17_47,N2_18_47,N2_19_47,N3_20_47,N3_21_48);
-- In matrix 2 adding FA to column 47 
	-- signal N3_22_47 : std_logic;
	-- signal N3_23_48 : std_logic;
	FA498 : full_adder port map (N2_20_47,N2_21_47,N2_22_47,N3_22_47,N3_23_48);
-- In matrix 2 adding FA to column 48 
	-- signal N3_0_48 : std_logic;
	-- signal N3_1_49 : std_logic;
	FA499 : full_adder port map (N0_38_48,N0_39_48,N0_40_48,N3_0_48,N3_1_49);
-- In matrix 2 adding FA to column 48 
	-- signal N3_2_48 : std_logic;
	-- signal N3_3_49 : std_logic;
	FA500 : full_adder port map (N0_41_48,N0_42_48,N0_43_48,N3_2_48,N3_3_49);
-- In matrix 2 adding FA to column 48 
	-- signal N3_4_48 : std_logic;
	-- signal N3_5_49 : std_logic;
	FA501 : full_adder port map (N0_44_48,N0_45_48,N0_46_48,N3_4_48,N3_5_49);
-- In matrix 2 adding FA to column 48 
	-- signal N3_6_48 : std_logic;
	-- signal N3_7_49 : std_logic;
	FA502 : full_adder port map (N0_47_48,N0_48_48,N2_0_48,N3_6_48,N3_7_49);
-- In matrix 2 adding FA to column 48 
	-- signal N3_8_48 : std_logic;
	-- signal N3_9_49 : std_logic;
	FA503 : full_adder port map (N2_1_48,N2_2_48,N2_3_48,N3_8_48,N3_9_49);
-- In matrix 2 adding FA to column 48 
	-- signal N3_10_48 : std_logic;
	-- signal N3_11_49 : std_logic;
	FA504 : full_adder port map (N2_4_48,N2_5_48,N2_6_48,N3_10_48,N3_11_49);
-- In matrix 2 adding FA to column 48 
	-- signal N3_12_48 : std_logic;
	-- signal N3_13_49 : std_logic;
	FA505 : full_adder port map (N2_7_48,N2_8_48,N2_9_48,N3_12_48,N3_13_49);
-- In matrix 2 adding FA to column 48 
	-- signal N3_14_48 : std_logic;
	-- signal N3_15_49 : std_logic;
	FA506 : full_adder port map (N2_10_48,N2_11_48,N2_12_48,N3_14_48,N3_15_49);
-- In matrix 2 adding FA to column 48 
	-- signal N3_16_48 : std_logic;
	-- signal N3_17_49 : std_logic;
	FA507 : full_adder port map (N2_13_48,N2_14_48,N2_15_48,N3_16_48,N3_17_49);
-- In matrix 2 adding FA to column 48 
	-- signal N3_18_48 : std_logic;
	-- signal N3_19_49 : std_logic;
	FA508 : full_adder port map (N2_16_48,N2_17_48,N2_18_48,N3_18_48,N3_19_49);
-- In matrix 2 adding FA to column 48 
	-- signal N3_20_48 : std_logic;
	-- signal N3_21_49 : std_logic;
	FA509 : full_adder port map (N2_19_48,N2_20_48,N2_21_48,N3_20_48,N3_21_49);
-- In matrix 2 adding FA to column 48 
	-- signal N3_22_48 : std_logic;
	-- signal N3_23_49 : std_logic;
	FA510 : full_adder port map (N2_22_48,N2_23_48,N2_24_48,N3_22_48,N3_23_49);
-- In matrix 2 adding FA to column 49 
	-- signal N3_0_49 : std_logic;
	-- signal N3_1_50 : std_logic;
	FA511 : full_adder port map (N0_41_49,N0_42_49,N0_43_49,N3_0_49,N3_1_50);
-- In matrix 2 adding FA to column 49 
	-- signal N3_2_49 : std_logic;
	-- signal N3_3_50 : std_logic;
	FA512 : full_adder port map (N0_44_49,N0_45_49,N0_46_49,N3_2_49,N3_3_50);
-- In matrix 2 adding FA to column 49 
	-- signal N3_4_49 : std_logic;
	-- signal N3_5_50 : std_logic;
	FA513 : full_adder port map (N0_47_49,N0_48_49,N0_49_49,N3_4_49,N3_5_50);
-- In matrix 2 adding FA to column 49 
	-- signal N3_6_49 : std_logic;
	-- signal N3_7_50 : std_logic;
	FA514 : full_adder port map (N2_0_49,N2_1_49,N2_2_49,N3_6_49,N3_7_50);
-- In matrix 2 adding FA to column 49 
	-- signal N3_8_49 : std_logic;
	-- signal N3_9_50 : std_logic;
	FA515 : full_adder port map (N2_3_49,N2_4_49,N2_5_49,N3_8_49,N3_9_50);
-- In matrix 2 adding FA to column 49 
	-- signal N3_10_49 : std_logic;
	-- signal N3_11_50 : std_logic;
	FA516 : full_adder port map (N2_6_49,N2_7_49,N2_8_49,N3_10_49,N3_11_50);
-- In matrix 2 adding FA to column 49 
	-- signal N3_12_49 : std_logic;
	-- signal N3_13_50 : std_logic;
	FA517 : full_adder port map (N2_9_49,N2_10_49,N2_11_49,N3_12_49,N3_13_50);
-- In matrix 2 adding FA to column 49 
	-- signal N3_14_49 : std_logic;
	-- signal N3_15_50 : std_logic;
	FA518 : full_adder port map (N2_12_49,N2_13_49,N2_14_49,N3_14_49,N3_15_50);
-- In matrix 2 adding FA to column 49 
	-- signal N3_16_49 : std_logic;
	-- signal N3_17_50 : std_logic;
	FA519 : full_adder port map (N2_15_49,N2_16_49,N2_17_49,N3_16_49,N3_17_50);
-- In matrix 2 adding FA to column 49 
	-- signal N3_18_49 : std_logic;
	-- signal N3_19_50 : std_logic;
	FA520 : full_adder port map (N2_18_49,N2_19_49,N2_20_49,N3_18_49,N3_19_50);
-- In matrix 2 adding FA to column 49 
	-- signal N3_20_49 : std_logic;
	-- signal N3_21_50 : std_logic;
	FA521 : full_adder port map (N2_21_49,N2_22_49,N2_23_49,N3_20_49,N3_21_50);
-- In matrix 2 adding FA to column 49 
	-- signal N3_22_49 : std_logic;
	-- signal N3_23_50 : std_logic;
	FA522 : full_adder port map (N2_24_49,N2_25_49,N2_26_49,N3_22_49,N3_23_50);
-- In matrix 2 adding FA to column 50 
	-- signal N3_0_50 : std_logic;
	-- signal N3_1_51 : std_logic;
	FA523 : full_adder port map (N0_44_50,N0_45_50,N0_46_50,N3_0_50,N3_1_51);
-- In matrix 2 adding FA to column 50 
	-- signal N3_2_50 : std_logic;
	-- signal N3_3_51 : std_logic;
	FA524 : full_adder port map (N0_47_50,N0_48_50,N0_49_50,N3_2_50,N3_3_51);
-- In matrix 2 adding FA to column 50 
	-- signal N3_4_50 : std_logic;
	-- signal N3_5_51 : std_logic;
	FA525 : full_adder port map (N0_50_50,N2_0_50,N2_1_50,N3_4_50,N3_5_51);
-- In matrix 2 adding FA to column 50 
	-- signal N3_6_50 : std_logic;
	-- signal N3_7_51 : std_logic;
	FA526 : full_adder port map (N2_2_50,N2_3_50,N2_4_50,N3_6_50,N3_7_51);
-- In matrix 2 adding FA to column 50 
	-- signal N3_8_50 : std_logic;
	-- signal N3_9_51 : std_logic;
	FA527 : full_adder port map (N2_5_50,N2_6_50,N2_7_50,N3_8_50,N3_9_51);
-- In matrix 2 adding FA to column 50 
	-- signal N3_10_50 : std_logic;
	-- signal N3_11_51 : std_logic;
	FA528 : full_adder port map (N2_8_50,N2_9_50,N2_10_50,N3_10_50,N3_11_51);
-- In matrix 2 adding FA to column 50 
	-- signal N3_12_50 : std_logic;
	-- signal N3_13_51 : std_logic;
	FA529 : full_adder port map (N2_11_50,N2_12_50,N2_13_50,N3_12_50,N3_13_51);
-- In matrix 2 adding FA to column 50 
	-- signal N3_14_50 : std_logic;
	-- signal N3_15_51 : std_logic;
	FA530 : full_adder port map (N2_14_50,N2_15_50,N2_16_50,N3_14_50,N3_15_51);
-- In matrix 2 adding FA to column 50 
	-- signal N3_16_50 : std_logic;
	-- signal N3_17_51 : std_logic;
	FA531 : full_adder port map (N2_17_50,N2_18_50,N2_19_50,N3_16_50,N3_17_51);
-- In matrix 2 adding FA to column 50 
	-- signal N3_18_50 : std_logic;
	-- signal N3_19_51 : std_logic;
	FA532 : full_adder port map (N2_20_50,N2_21_50,N2_22_50,N3_18_50,N3_19_51);
-- In matrix 2 adding FA to column 50 
	-- signal N3_20_50 : std_logic;
	-- signal N3_21_51 : std_logic;
	FA533 : full_adder port map (N2_23_50,N2_24_50,N2_25_50,N3_20_50,N3_21_51);
-- In matrix 2 adding FA to column 50 
	-- signal N3_22_50 : std_logic;
	-- signal N3_23_51 : std_logic;
	FA534 : full_adder port map (N2_26_50,N2_27_50,N2_28_50,N3_22_50,N3_23_51);
-- In matrix 2 adding FA to column 51 
	-- signal N3_0_51 : std_logic;
	-- signal N3_1_52 : std_logic;
	FA535 : full_adder port map (N0_47_51,N0_48_51,N0_49_51,N3_0_51,N3_1_52);
-- In matrix 2 adding FA to column 51 
	-- signal N3_2_51 : std_logic;
	-- signal N3_3_52 : std_logic;
	FA536 : full_adder port map (N0_50_51,N0_51_51,N2_0_51,N3_2_51,N3_3_52);
-- In matrix 2 adding FA to column 51 
	-- signal N3_4_51 : std_logic;
	-- signal N3_5_52 : std_logic;
	FA537 : full_adder port map (N2_1_51,N2_2_51,N2_3_51,N3_4_51,N3_5_52);
-- In matrix 2 adding FA to column 51 
	-- signal N3_6_51 : std_logic;
	-- signal N3_7_52 : std_logic;
	FA538 : full_adder port map (N2_4_51,N2_5_51,N2_6_51,N3_6_51,N3_7_52);
-- In matrix 2 adding FA to column 51 
	-- signal N3_8_51 : std_logic;
	-- signal N3_9_52 : std_logic;
	FA539 : full_adder port map (N2_7_51,N2_8_51,N2_9_51,N3_8_51,N3_9_52);
-- In matrix 2 adding FA to column 51 
	-- signal N3_10_51 : std_logic;
	-- signal N3_11_52 : std_logic;
	FA540 : full_adder port map (N2_10_51,N2_11_51,N2_12_51,N3_10_51,N3_11_52);
-- In matrix 2 adding FA to column 51 
	-- signal N3_12_51 : std_logic;
	-- signal N3_13_52 : std_logic;
	FA541 : full_adder port map (N2_13_51,N2_14_51,N2_15_51,N3_12_51,N3_13_52);
-- In matrix 2 adding FA to column 51 
	-- signal N3_14_51 : std_logic;
	-- signal N3_15_52 : std_logic;
	FA542 : full_adder port map (N2_16_51,N2_17_51,N2_18_51,N3_14_51,N3_15_52);
-- In matrix 2 adding FA to column 51 
	-- signal N3_16_51 : std_logic;
	-- signal N3_17_52 : std_logic;
	FA543 : full_adder port map (N2_19_51,N2_20_51,N2_21_51,N3_16_51,N3_17_52);
-- In matrix 2 adding FA to column 51 
	-- signal N3_18_51 : std_logic;
	-- signal N3_19_52 : std_logic;
	FA544 : full_adder port map (N2_22_51,N2_23_51,N2_24_51,N3_18_51,N3_19_52);
-- In matrix 2 adding FA to column 51 
	-- signal N3_20_51 : std_logic;
	-- signal N3_21_52 : std_logic;
	FA545 : full_adder port map (N2_25_51,N2_26_51,N2_27_51,N3_20_51,N3_21_52);
-- In matrix 2 adding FA to column 51 
	-- signal N3_22_51 : std_logic;
	-- signal N3_23_52 : std_logic;
	FA546 : full_adder port map (N2_28_51,N2_29_51,N2_30_51,N3_22_51,N3_23_52);
-- In matrix 2 adding FA to column 52 
	-- signal N3_0_52 : std_logic;
	-- signal N3_1_53 : std_logic;
	FA547 : full_adder port map (N0_50_52,N0_51_52,N0_52_52,N3_0_52,N3_1_53);
-- In matrix 2 adding FA to column 52 
	-- signal N3_2_52 : std_logic;
	-- signal N3_3_53 : std_logic;
	FA548 : full_adder port map (N2_0_52,N2_1_52,N2_2_52,N3_2_52,N3_3_53);
-- In matrix 2 adding FA to column 52 
	-- signal N3_4_52 : std_logic;
	-- signal N3_5_53 : std_logic;
	FA549 : full_adder port map (N2_3_52,N2_4_52,N2_5_52,N3_4_52,N3_5_53);
-- In matrix 2 adding FA to column 52 
	-- signal N3_6_52 : std_logic;
	-- signal N3_7_53 : std_logic;
	FA550 : full_adder port map (N2_6_52,N2_7_52,N2_8_52,N3_6_52,N3_7_53);
-- In matrix 2 adding FA to column 52 
	-- signal N3_8_52 : std_logic;
	-- signal N3_9_53 : std_logic;
	FA551 : full_adder port map (N2_9_52,N2_10_52,N2_11_52,N3_8_52,N3_9_53);
-- In matrix 2 adding FA to column 52 
	-- signal N3_10_52 : std_logic;
	-- signal N3_11_53 : std_logic;
	FA552 : full_adder port map (N2_12_52,N2_13_52,N2_14_52,N3_10_52,N3_11_53);
-- In matrix 2 adding FA to column 52 
	-- signal N3_12_52 : std_logic;
	-- signal N3_13_53 : std_logic;
	FA553 : full_adder port map (N2_15_52,N2_16_52,N2_17_52,N3_12_52,N3_13_53);
-- In matrix 2 adding FA to column 52 
	-- signal N3_14_52 : std_logic;
	-- signal N3_15_53 : std_logic;
	FA554 : full_adder port map (N2_18_52,N2_19_52,N2_20_52,N3_14_52,N3_15_53);
-- In matrix 2 adding FA to column 52 
	-- signal N3_16_52 : std_logic;
	-- signal N3_17_53 : std_logic;
	FA555 : full_adder port map (N2_21_52,N2_22_52,N2_23_52,N3_16_52,N3_17_53);
-- In matrix 2 adding FA to column 52 
	-- signal N3_18_52 : std_logic;
	-- signal N3_19_53 : std_logic;
	FA556 : full_adder port map (N2_24_52,N2_25_52,N2_26_52,N3_18_52,N3_19_53);
-- In matrix 2 adding FA to column 52 
	-- signal N3_20_52 : std_logic;
	-- signal N3_21_53 : std_logic;
	FA557 : full_adder port map (N2_27_52,N2_28_52,N2_29_52,N3_20_52,N3_21_53);
-- In matrix 2 adding FA to column 52 
	-- signal N3_22_52 : std_logic;
	-- signal N3_23_53 : std_logic;
	FA558 : full_adder port map (N2_30_52,N2_31_52,N2_32_52,N3_22_52,N3_23_53);
-- In matrix 2 adding FA to column 53 
	-- signal N3_0_53 : std_logic;
	-- signal N3_1_54 : std_logic;
	FA559 : full_adder port map (N0_51_53,N0_52_53,N2_0_53,N3_0_53,N3_1_54);
-- In matrix 2 adding FA to column 53 
	-- signal N3_2_53 : std_logic;
	-- signal N3_3_54 : std_logic;
	FA560 : full_adder port map (N2_1_53,N2_2_53,N2_3_53,N3_2_53,N3_3_54);
-- In matrix 2 adding FA to column 53 
	-- signal N3_4_53 : std_logic;
	-- signal N3_5_54 : std_logic;
	FA561 : full_adder port map (N2_4_53,N2_5_53,N2_6_53,N3_4_53,N3_5_54);
-- In matrix 2 adding FA to column 53 
	-- signal N3_6_53 : std_logic;
	-- signal N3_7_54 : std_logic;
	FA562 : full_adder port map (N2_7_53,N2_8_53,N2_9_53,N3_6_53,N3_7_54);
-- In matrix 2 adding FA to column 53 
	-- signal N3_8_53 : std_logic;
	-- signal N3_9_54 : std_logic;
	FA563 : full_adder port map (N2_10_53,N2_11_53,N2_12_53,N3_8_53,N3_9_54);
-- In matrix 2 adding FA to column 53 
	-- signal N3_10_53 : std_logic;
	-- signal N3_11_54 : std_logic;
	FA564 : full_adder port map (N2_13_53,N2_14_53,N2_15_53,N3_10_53,N3_11_54);
-- In matrix 2 adding FA to column 53 
	-- signal N3_12_53 : std_logic;
	-- signal N3_13_54 : std_logic;
	FA565 : full_adder port map (N2_16_53,N2_17_53,N2_18_53,N3_12_53,N3_13_54);
-- In matrix 2 adding FA to column 53 
	-- signal N3_14_53 : std_logic;
	-- signal N3_15_54 : std_logic;
	FA566 : full_adder port map (N2_19_53,N2_20_53,N2_21_53,N3_14_53,N3_15_54);
-- In matrix 2 adding FA to column 53 
	-- signal N3_16_53 : std_logic;
	-- signal N3_17_54 : std_logic;
	FA567 : full_adder port map (N2_22_53,N2_23_53,N2_24_53,N3_16_53,N3_17_54);
-- In matrix 2 adding FA to column 53 
	-- signal N3_18_53 : std_logic;
	-- signal N3_19_54 : std_logic;
	FA568 : full_adder port map (N2_25_53,N2_26_53,N2_27_53,N3_18_53,N3_19_54);
-- In matrix 2 adding FA to column 53 
	-- signal N3_20_53 : std_logic;
	-- signal N3_21_54 : std_logic;
	FA569 : full_adder port map (N2_28_53,N2_29_53,N2_30_53,N3_20_53,N3_21_54);
-- In matrix 2 adding FA to column 53 
	-- signal N3_22_53 : std_logic;
	-- signal N3_23_54 : std_logic;
	FA570 : full_adder port map (N2_31_53,N2_32_53,N2_33_53,N3_22_53,N3_23_54);
-- In matrix 2 adding FA to column 54 
	-- signal N3_0_54 : std_logic;
	-- signal N3_1_55 : std_logic;
	FA571 : full_adder port map (N0_50_54,N0_51_54,N0_52_54,N3_0_54,N3_1_55);
-- In matrix 2 adding FA to column 54 
	-- signal N3_2_54 : std_logic;
	-- signal N3_3_55 : std_logic;
	FA572 : full_adder port map (N2_0_54,N2_1_54,N2_2_54,N3_2_54,N3_3_55);
-- In matrix 2 adding FA to column 54 
	-- signal N3_4_54 : std_logic;
	-- signal N3_5_55 : std_logic;
	FA573 : full_adder port map (N2_3_54,N2_4_54,N2_5_54,N3_4_54,N3_5_55);
-- In matrix 2 adding FA to column 54 
	-- signal N3_6_54 : std_logic;
	-- signal N3_7_55 : std_logic;
	FA574 : full_adder port map (N2_6_54,N2_7_54,N2_8_54,N3_6_54,N3_7_55);
-- In matrix 2 adding FA to column 54 
	-- signal N3_8_54 : std_logic;
	-- signal N3_9_55 : std_logic;
	FA575 : full_adder port map (N2_9_54,N2_10_54,N2_11_54,N3_8_54,N3_9_55);
-- In matrix 2 adding FA to column 54 
	-- signal N3_10_54 : std_logic;
	-- signal N3_11_55 : std_logic;
	FA576 : full_adder port map (N2_12_54,N2_13_54,N2_14_54,N3_10_54,N3_11_55);
-- In matrix 2 adding FA to column 54 
	-- signal N3_12_54 : std_logic;
	-- signal N3_13_55 : std_logic;
	FA577 : full_adder port map (N2_15_54,N2_16_54,N2_17_54,N3_12_54,N3_13_55);
-- In matrix 2 adding FA to column 54 
	-- signal N3_14_54 : std_logic;
	-- signal N3_15_55 : std_logic;
	FA578 : full_adder port map (N2_18_54,N2_19_54,N2_20_54,N3_14_54,N3_15_55);
-- In matrix 2 adding FA to column 54 
	-- signal N3_16_54 : std_logic;
	-- signal N3_17_55 : std_logic;
	FA579 : full_adder port map (N2_21_54,N2_22_54,N2_23_54,N3_16_54,N3_17_55);
-- In matrix 2 adding FA to column 54 
	-- signal N3_18_54 : std_logic;
	-- signal N3_19_55 : std_logic;
	FA580 : full_adder port map (N2_24_54,N2_25_54,N2_26_54,N3_18_54,N3_19_55);
-- In matrix 2 adding FA to column 54 
	-- signal N3_20_54 : std_logic;
	-- signal N3_21_55 : std_logic;
	FA581 : full_adder port map (N2_27_54,N2_28_54,N2_29_54,N3_20_54,N3_21_55);
-- In matrix 2 adding FA to column 54 
	-- signal N3_22_54 : std_logic;
	-- signal N3_23_55 : std_logic;
	FA582 : full_adder port map (N2_30_54,N2_31_54,N2_33_54,N3_22_54,N3_23_55);
-- In matrix 2 adding FA to column 55 
	-- signal N3_0_55 : std_logic;
	-- signal N3_1_56 : std_logic;
	FA583 : full_adder port map (N0_48_55,N0_49_55,N0_50_55,N3_0_55,N3_1_56);
-- In matrix 2 adding FA to column 55 
	-- signal N3_2_55 : std_logic;
	-- signal N3_3_56 : std_logic;
	FA584 : full_adder port map (N0_51_55,N0_52_55,N2_0_55,N3_2_55,N3_3_56);
-- In matrix 2 adding FA to column 55 
	-- signal N3_4_55 : std_logic;
	-- signal N3_5_56 : std_logic;
	FA585 : full_adder port map (N2_1_55,N2_2_55,N2_3_55,N3_4_55,N3_5_56);
-- In matrix 2 adding FA to column 55 
	-- signal N3_6_55 : std_logic;
	-- signal N3_7_56 : std_logic;
	FA586 : full_adder port map (N2_4_55,N2_5_55,N2_6_55,N3_6_55,N3_7_56);
-- In matrix 2 adding FA to column 55 
	-- signal N3_8_55 : std_logic;
	-- signal N3_9_56 : std_logic;
	FA587 : full_adder port map (N2_7_55,N2_8_55,N2_9_55,N3_8_55,N3_9_56);
-- In matrix 2 adding FA to column 55 
	-- signal N3_10_55 : std_logic;
	-- signal N3_11_56 : std_logic;
	FA588 : full_adder port map (N2_10_55,N2_11_55,N2_12_55,N3_10_55,N3_11_56);
-- In matrix 2 adding FA to column 55 
	-- signal N3_12_55 : std_logic;
	-- signal N3_13_56 : std_logic;
	FA589 : full_adder port map (N2_13_55,N2_14_55,N2_15_55,N3_12_55,N3_13_56);
-- In matrix 2 adding FA to column 55 
	-- signal N3_14_55 : std_logic;
	-- signal N3_15_56 : std_logic;
	FA590 : full_adder port map (N2_16_55,N2_17_55,N2_18_55,N3_14_55,N3_15_56);
-- In matrix 2 adding FA to column 55 
	-- signal N3_16_55 : std_logic;
	-- signal N3_17_56 : std_logic;
	FA591 : full_adder port map (N2_19_55,N2_20_55,N2_21_55,N3_16_55,N3_17_56);
-- In matrix 2 adding FA to column 55 
	-- signal N3_18_55 : std_logic;
	-- signal N3_19_56 : std_logic;
	FA592 : full_adder port map (N2_22_55,N2_23_55,N2_24_55,N3_18_55,N3_19_56);
-- In matrix 2 adding FA to column 55 
	-- signal N3_20_55 : std_logic;
	-- signal N3_21_56 : std_logic;
	FA593 : full_adder port map (N2_25_55,N2_26_55,N2_27_55,N3_20_55,N3_21_56);
-- In matrix 2 adding FA to column 55 
	-- signal N3_22_55 : std_logic;
	-- signal N3_23_56 : std_logic;
	FA594 : full_adder port map (N2_28_55,N2_29_55,N2_31_55,N3_22_55,N3_23_56);
-- In matrix 2 adding FA to column 56 
	-- signal N3_0_56 : std_logic;
	-- signal N3_1_57 : std_logic;
	FA595 : full_adder port map (N0_46_56,N0_47_56,N0_48_56,N3_0_56,N3_1_57);
-- In matrix 2 adding FA to column 56 
	-- signal N3_2_56 : std_logic;
	-- signal N3_3_57 : std_logic;
	FA596 : full_adder port map (N0_49_56,N0_50_56,N0_51_56,N3_2_56,N3_3_57);
-- In matrix 2 adding FA to column 56 
	-- signal N3_4_56 : std_logic;
	-- signal N3_5_57 : std_logic;
	FA597 : full_adder port map (N0_52_56,N2_0_56,N2_1_56,N3_4_56,N3_5_57);
-- In matrix 2 adding FA to column 56 
	-- signal N3_6_56 : std_logic;
	-- signal N3_7_57 : std_logic;
	FA598 : full_adder port map (N2_2_56,N2_3_56,N2_4_56,N3_6_56,N3_7_57);
-- In matrix 2 adding FA to column 56 
	-- signal N3_8_56 : std_logic;
	-- signal N3_9_57 : std_logic;
	FA599 : full_adder port map (N2_5_56,N2_6_56,N2_7_56,N3_8_56,N3_9_57);
-- In matrix 2 adding FA to column 56 
	-- signal N3_10_56 : std_logic;
	-- signal N3_11_57 : std_logic;
	FA600 : full_adder port map (N2_8_56,N2_9_56,N2_10_56,N3_10_56,N3_11_57);
-- In matrix 2 adding FA to column 56 
	-- signal N3_12_56 : std_logic;
	-- signal N3_13_57 : std_logic;
	FA601 : full_adder port map (N2_11_56,N2_12_56,N2_13_56,N3_12_56,N3_13_57);
-- In matrix 2 adding FA to column 56 
	-- signal N3_14_56 : std_logic;
	-- signal N3_15_57 : std_logic;
	FA602 : full_adder port map (N2_14_56,N2_15_56,N2_16_56,N3_14_56,N3_15_57);
-- In matrix 2 adding FA to column 56 
	-- signal N3_16_56 : std_logic;
	-- signal N3_17_57 : std_logic;
	FA603 : full_adder port map (N2_17_56,N2_18_56,N2_19_56,N3_16_56,N3_17_57);
-- In matrix 2 adding FA to column 56 
	-- signal N3_18_56 : std_logic;
	-- signal N3_19_57 : std_logic;
	FA604 : full_adder port map (N2_20_56,N2_21_56,N2_22_56,N3_18_56,N3_19_57);
-- In matrix 2 adding FA to column 56 
	-- signal N3_20_56 : std_logic;
	-- signal N3_21_57 : std_logic;
	FA605 : full_adder port map (N2_23_56,N2_24_56,N2_25_56,N3_20_56,N3_21_57);
-- In matrix 2 adding FA to column 56 
	-- signal N3_22_56 : std_logic;
	-- signal N3_23_57 : std_logic;
	FA606 : full_adder port map (N2_26_56,N2_27_56,N2_29_56,N3_22_56,N3_23_57);
-- In matrix 2 adding FA to column 57 
	-- signal N3_0_57 : std_logic;
	-- signal N3_1_58 : std_logic;
	FA607 : full_adder port map (N0_44_57,N0_45_57,N0_46_57,N3_0_57,N3_1_58);
-- In matrix 2 adding FA to column 57 
	-- signal N3_2_57 : std_logic;
	-- signal N3_3_58 : std_logic;
	FA608 : full_adder port map (N0_47_57,N0_48_57,N0_49_57,N3_2_57,N3_3_58);
-- In matrix 2 adding FA to column 57 
	-- signal N3_4_57 : std_logic;
	-- signal N3_5_58 : std_logic;
	FA609 : full_adder port map (N0_50_57,N0_51_57,N0_52_57,N3_4_57,N3_5_58);
-- In matrix 2 adding FA to column 57 
	-- signal N3_6_57 : std_logic;
	-- signal N3_7_58 : std_logic;
	FA610 : full_adder port map (N2_0_57,N2_1_57,N2_2_57,N3_6_57,N3_7_58);
-- In matrix 2 adding FA to column 57 
	-- signal N3_8_57 : std_logic;
	-- signal N3_9_58 : std_logic;
	FA611 : full_adder port map (N2_3_57,N2_4_57,N2_5_57,N3_8_57,N3_9_58);
-- In matrix 2 adding FA to column 57 
	-- signal N3_10_57 : std_logic;
	-- signal N3_11_58 : std_logic;
	FA612 : full_adder port map (N2_6_57,N2_7_57,N2_8_57,N3_10_57,N3_11_58);
-- In matrix 2 adding FA to column 57 
	-- signal N3_12_57 : std_logic;
	-- signal N3_13_58 : std_logic;
	FA613 : full_adder port map (N2_9_57,N2_10_57,N2_11_57,N3_12_57,N3_13_58);
-- In matrix 2 adding FA to column 57 
	-- signal N3_14_57 : std_logic;
	-- signal N3_15_58 : std_logic;
	FA614 : full_adder port map (N2_12_57,N2_13_57,N2_14_57,N3_14_57,N3_15_58);
-- In matrix 2 adding FA to column 57 
	-- signal N3_16_57 : std_logic;
	-- signal N3_17_58 : std_logic;
	FA615 : full_adder port map (N2_15_57,N2_16_57,N2_17_57,N3_16_57,N3_17_58);
-- In matrix 2 adding FA to column 57 
	-- signal N3_18_57 : std_logic;
	-- signal N3_19_58 : std_logic;
	FA616 : full_adder port map (N2_18_57,N2_19_57,N2_20_57,N3_18_57,N3_19_58);
-- In matrix 2 adding FA to column 57 
	-- signal N3_20_57 : std_logic;
	-- signal N3_21_58 : std_logic;
	FA617 : full_adder port map (N2_21_57,N2_22_57,N2_23_57,N3_20_57,N3_21_58);
-- In matrix 2 adding FA to column 57 
	-- signal N3_22_57 : std_logic;
	-- signal N3_23_58 : std_logic;
	FA618 : full_adder port map (N2_24_57,N2_25_57,N2_27_57,N3_22_57,N3_23_58);
-- In matrix 2 adding FA to column 58 
	-- signal N3_0_58 : std_logic;
	-- signal N3_1_59 : std_logic;
	FA619 : full_adder port map (N0_42_58,N0_43_58,N0_44_58,N3_0_58,N3_1_59);
-- In matrix 2 adding FA to column 58 
	-- signal N3_2_58 : std_logic;
	-- signal N3_3_59 : std_logic;
	FA620 : full_adder port map (N0_45_58,N0_46_58,N0_47_58,N3_2_58,N3_3_59);
-- In matrix 2 adding FA to column 58 
	-- signal N3_4_58 : std_logic;
	-- signal N3_5_59 : std_logic;
	FA621 : full_adder port map (N0_48_58,N0_49_58,N0_50_58,N3_4_58,N3_5_59);
-- In matrix 2 adding FA to column 58 
	-- signal N3_6_58 : std_logic;
	-- signal N3_7_59 : std_logic;
	FA622 : full_adder port map (N0_51_58,N0_52_58,N2_0_58,N3_6_58,N3_7_59);
-- In matrix 2 adding FA to column 58 
	-- signal N3_8_58 : std_logic;
	-- signal N3_9_59 : std_logic;
	FA623 : full_adder port map (N2_1_58,N2_2_58,N2_3_58,N3_8_58,N3_9_59);
-- In matrix 2 adding FA to column 58 
	-- signal N3_10_58 : std_logic;
	-- signal N3_11_59 : std_logic;
	FA624 : full_adder port map (N2_4_58,N2_5_58,N2_6_58,N3_10_58,N3_11_59);
-- In matrix 2 adding FA to column 58 
	-- signal N3_12_58 : std_logic;
	-- signal N3_13_59 : std_logic;
	FA625 : full_adder port map (N2_7_58,N2_8_58,N2_9_58,N3_12_58,N3_13_59);
-- In matrix 2 adding FA to column 58 
	-- signal N3_14_58 : std_logic;
	-- signal N3_15_59 : std_logic;
	FA626 : full_adder port map (N2_10_58,N2_11_58,N2_12_58,N3_14_58,N3_15_59);
-- In matrix 2 adding FA to column 58 
	-- signal N3_16_58 : std_logic;
	-- signal N3_17_59 : std_logic;
	FA627 : full_adder port map (N2_13_58,N2_14_58,N2_15_58,N3_16_58,N3_17_59);
-- In matrix 2 adding FA to column 58 
	-- signal N3_18_58 : std_logic;
	-- signal N3_19_59 : std_logic;
	FA628 : full_adder port map (N2_16_58,N2_17_58,N2_18_58,N3_18_58,N3_19_59);
-- In matrix 2 adding FA to column 58 
	-- signal N3_20_58 : std_logic;
	-- signal N3_21_59 : std_logic;
	FA629 : full_adder port map (N2_19_58,N2_20_58,N2_21_58,N3_20_58,N3_21_59);
-- In matrix 2 adding FA to column 58 
	-- signal N3_22_58 : std_logic;
	-- signal N3_23_59 : std_logic;
	FA630 : full_adder port map (N2_22_58,N2_23_58,N2_25_58,N3_22_58,N3_23_59);
-- In matrix 2 adding FA to column 59 
	-- signal N3_0_59 : std_logic;
	-- signal N3_1_60 : std_logic;
	FA631 : full_adder port map (N0_40_59,N0_41_59,N0_42_59,N3_0_59,N3_1_60);
-- In matrix 2 adding FA to column 59 
	-- signal N3_2_59 : std_logic;
	-- signal N3_3_60 : std_logic;
	FA632 : full_adder port map (N0_43_59,N0_44_59,N0_45_59,N3_2_59,N3_3_60);
-- In matrix 2 adding FA to column 59 
	-- signal N3_4_59 : std_logic;
	-- signal N3_5_60 : std_logic;
	FA633 : full_adder port map (N0_46_59,N0_47_59,N0_48_59,N3_4_59,N3_5_60);
-- In matrix 2 adding FA to column 59 
	-- signal N3_6_59 : std_logic;
	-- signal N3_7_60 : std_logic;
	FA634 : full_adder port map (N0_49_59,N0_50_59,N0_51_59,N3_6_59,N3_7_60);
-- In matrix 2 adding FA to column 59 
	-- signal N3_8_59 : std_logic;
	-- signal N3_9_60 : std_logic;
	FA635 : full_adder port map (N0_52_59,N2_0_59,N2_1_59,N3_8_59,N3_9_60);
-- In matrix 2 adding FA to column 59 
	-- signal N3_10_59 : std_logic;
	-- signal N3_11_60 : std_logic;
	FA636 : full_adder port map (N2_2_59,N2_3_59,N2_4_59,N3_10_59,N3_11_60);
-- In matrix 2 adding FA to column 59 
	-- signal N3_12_59 : std_logic;
	-- signal N3_13_60 : std_logic;
	FA637 : full_adder port map (N2_5_59,N2_6_59,N2_7_59,N3_12_59,N3_13_60);
-- In matrix 2 adding FA to column 59 
	-- signal N3_14_59 : std_logic;
	-- signal N3_15_60 : std_logic;
	FA638 : full_adder port map (N2_8_59,N2_9_59,N2_10_59,N3_14_59,N3_15_60);
-- In matrix 2 adding FA to column 59 
	-- signal N3_16_59 : std_logic;
	-- signal N3_17_60 : std_logic;
	FA639 : full_adder port map (N2_11_59,N2_12_59,N2_13_59,N3_16_59,N3_17_60);
-- In matrix 2 adding FA to column 59 
	-- signal N3_18_59 : std_logic;
	-- signal N3_19_60 : std_logic;
	FA640 : full_adder port map (N2_14_59,N2_15_59,N2_16_59,N3_18_59,N3_19_60);
-- In matrix 2 adding FA to column 59 
	-- signal N3_20_59 : std_logic;
	-- signal N3_21_60 : std_logic;
	FA641 : full_adder port map (N2_17_59,N2_18_59,N2_19_59,N3_20_59,N3_21_60);
-- In matrix 2 adding FA to column 59 
	-- signal N3_22_59 : std_logic;
	-- signal N3_23_60 : std_logic;
	FA642 : full_adder port map (N2_20_59,N2_21_59,N2_23_59,N3_22_59,N3_23_60);
-- In matrix 2 adding FA to column 60 
	-- signal N3_0_60 : std_logic;
	-- signal N3_1_61 : std_logic;
	FA643 : full_adder port map (N0_38_60,N0_39_60,N0_40_60,N3_0_60,N3_1_61);
-- In matrix 2 adding FA to column 60 
	-- signal N3_2_60 : std_logic;
	-- signal N3_3_61 : std_logic;
	FA644 : full_adder port map (N0_41_60,N0_42_60,N0_43_60,N3_2_60,N3_3_61);
-- In matrix 2 adding FA to column 60 
	-- signal N3_4_60 : std_logic;
	-- signal N3_5_61 : std_logic;
	FA645 : full_adder port map (N0_44_60,N0_45_60,N0_46_60,N3_4_60,N3_5_61);
-- In matrix 2 adding FA to column 60 
	-- signal N3_6_60 : std_logic;
	-- signal N3_7_61 : std_logic;
	FA646 : full_adder port map (N0_47_60,N0_48_60,N0_49_60,N3_6_60,N3_7_61);
-- In matrix 2 adding FA to column 60 
	-- signal N3_8_60 : std_logic;
	-- signal N3_9_61 : std_logic;
	FA647 : full_adder port map (N0_50_60,N0_51_60,N0_52_60,N3_8_60,N3_9_61);
-- In matrix 2 adding FA to column 60 
	-- signal N3_10_60 : std_logic;
	-- signal N3_11_61 : std_logic;
	FA648 : full_adder port map (N2_0_60,N2_1_60,N2_2_60,N3_10_60,N3_11_61);
-- In matrix 2 adding FA to column 60 
	-- signal N3_12_60 : std_logic;
	-- signal N3_13_61 : std_logic;
	FA649 : full_adder port map (N2_3_60,N2_4_60,N2_5_60,N3_12_60,N3_13_61);
-- In matrix 2 adding FA to column 60 
	-- signal N3_14_60 : std_logic;
	-- signal N3_15_61 : std_logic;
	FA650 : full_adder port map (N2_6_60,N2_7_60,N2_8_60,N3_14_60,N3_15_61);
-- In matrix 2 adding FA to column 60 
	-- signal N3_16_60 : std_logic;
	-- signal N3_17_61 : std_logic;
	FA651 : full_adder port map (N2_9_60,N2_10_60,N2_11_60,N3_16_60,N3_17_61);
-- In matrix 2 adding FA to column 60 
	-- signal N3_18_60 : std_logic;
	-- signal N3_19_61 : std_logic;
	FA652 : full_adder port map (N2_12_60,N2_13_60,N2_14_60,N3_18_60,N3_19_61);
-- In matrix 2 adding FA to column 60 
	-- signal N3_20_60 : std_logic;
	-- signal N3_21_61 : std_logic;
	FA653 : full_adder port map (N2_15_60,N2_16_60,N2_17_60,N3_20_60,N3_21_61);
-- In matrix 2 adding FA to column 60 
	-- signal N3_22_60 : std_logic;
	-- signal N3_23_61 : std_logic;
	FA654 : full_adder port map (N2_18_60,N2_19_60,N2_21_60,N3_22_60,N3_23_61);
-- In matrix 2 adding FA to column 61 
	-- signal N3_0_61 : std_logic;
	-- signal N3_1_62 : std_logic;
	FA655 : full_adder port map (N0_36_61,N0_37_61,N0_38_61,N3_0_61,N3_1_62);
-- In matrix 2 adding FA to column 61 
	-- signal N3_2_61 : std_logic;
	-- signal N3_3_62 : std_logic;
	FA656 : full_adder port map (N0_39_61,N0_40_61,N0_41_61,N3_2_61,N3_3_62);
-- In matrix 2 adding FA to column 61 
	-- signal N3_4_61 : std_logic;
	-- signal N3_5_62 : std_logic;
	FA657 : full_adder port map (N0_42_61,N0_43_61,N0_44_61,N3_4_61,N3_5_62);
-- In matrix 2 adding FA to column 61 
	-- signal N3_6_61 : std_logic;
	-- signal N3_7_62 : std_logic;
	FA658 : full_adder port map (N0_45_61,N0_46_61,N0_47_61,N3_6_61,N3_7_62);
-- In matrix 2 adding FA to column 61 
	-- signal N3_8_61 : std_logic;
	-- signal N3_9_62 : std_logic;
	FA659 : full_adder port map (N0_48_61,N0_49_61,N0_50_61,N3_8_61,N3_9_62);
-- In matrix 2 adding FA to column 61 
	-- signal N3_10_61 : std_logic;
	-- signal N3_11_62 : std_logic;
	FA660 : full_adder port map (N0_51_61,N0_52_61,N2_0_61,N3_10_61,N3_11_62);
-- In matrix 2 adding FA to column 61 
	-- signal N3_12_61 : std_logic;
	-- signal N3_13_62 : std_logic;
	FA661 : full_adder port map (N2_1_61,N2_2_61,N2_3_61,N3_12_61,N3_13_62);
-- In matrix 2 adding FA to column 61 
	-- signal N3_14_61 : std_logic;
	-- signal N3_15_62 : std_logic;
	FA662 : full_adder port map (N2_4_61,N2_5_61,N2_6_61,N3_14_61,N3_15_62);
-- In matrix 2 adding FA to column 61 
	-- signal N3_16_61 : std_logic;
	-- signal N3_17_62 : std_logic;
	FA663 : full_adder port map (N2_7_61,N2_8_61,N2_9_61,N3_16_61,N3_17_62);
-- In matrix 2 adding FA to column 61 
	-- signal N3_18_61 : std_logic;
	-- signal N3_19_62 : std_logic;
	FA664 : full_adder port map (N2_10_61,N2_11_61,N2_12_61,N3_18_61,N3_19_62);
-- In matrix 2 adding FA to column 61 
	-- signal N3_20_61 : std_logic;
	-- signal N3_21_62 : std_logic;
	FA665 : full_adder port map (N2_13_61,N2_14_61,N2_15_61,N3_20_61,N3_21_62);
-- In matrix 2 adding FA to column 61 
	-- signal N3_22_61 : std_logic;
	-- signal N3_23_62 : std_logic;
	FA666 : full_adder port map (N2_16_61,N2_17_61,N2_19_61,N3_22_61,N3_23_62);
-- In matrix 2 adding FA to column 62 
	-- signal N3_0_62 : std_logic;
	-- signal N3_1_63 : std_logic;
	FA667 : full_adder port map (N0_34_62,N0_35_62,N0_36_62,N3_0_62,N3_1_63);
-- In matrix 2 adding FA to column 62 
	-- signal N3_2_62 : std_logic;
	-- signal N3_3_63 : std_logic;
	FA668 : full_adder port map (N0_37_62,N0_38_62,N0_39_62,N3_2_62,N3_3_63);
-- In matrix 2 adding FA to column 62 
	-- signal N3_4_62 : std_logic;
	-- signal N3_5_63 : std_logic;
	FA669 : full_adder port map (N0_40_62,N0_41_62,N0_42_62,N3_4_62,N3_5_63);
-- In matrix 2 adding FA to column 62 
	-- signal N3_6_62 : std_logic;
	-- signal N3_7_63 : std_logic;
	FA670 : full_adder port map (N0_43_62,N0_44_62,N0_45_62,N3_6_62,N3_7_63);
-- In matrix 2 adding FA to column 62 
	-- signal N3_8_62 : std_logic;
	-- signal N3_9_63 : std_logic;
	FA671 : full_adder port map (N0_46_62,N0_47_62,N0_48_62,N3_8_62,N3_9_63);
-- In matrix 2 adding FA to column 62 
	-- signal N3_10_62 : std_logic;
	-- signal N3_11_63 : std_logic;
	FA672 : full_adder port map (N0_49_62,N0_50_62,N0_51_62,N3_10_62,N3_11_63);
-- In matrix 2 adding FA to column 62 
	-- signal N3_12_62 : std_logic;
	-- signal N3_13_63 : std_logic;
	FA673 : full_adder port map (N0_52_62,N2_0_62,N2_1_62,N3_12_62,N3_13_63);
-- In matrix 2 adding FA to column 62 
	-- signal N3_14_62 : std_logic;
	-- signal N3_15_63 : std_logic;
	FA674 : full_adder port map (N2_2_62,N2_3_62,N2_4_62,N3_14_62,N3_15_63);
-- In matrix 2 adding FA to column 62 
	-- signal N3_16_62 : std_logic;
	-- signal N3_17_63 : std_logic;
	FA675 : full_adder port map (N2_5_62,N2_6_62,N2_7_62,N3_16_62,N3_17_63);
-- In matrix 2 adding FA to column 62 
	-- signal N3_18_62 : std_logic;
	-- signal N3_19_63 : std_logic;
	FA676 : full_adder port map (N2_8_62,N2_9_62,N2_10_62,N3_18_62,N3_19_63);
-- In matrix 2 adding FA to column 62 
	-- signal N3_20_62 : std_logic;
	-- signal N3_21_63 : std_logic;
	FA677 : full_adder port map (N2_11_62,N2_12_62,N2_13_62,N3_20_62,N3_21_63);
-- In matrix 2 adding FA to column 62 
	-- signal N3_22_62 : std_logic;
	-- signal N3_23_63 : std_logic;
	FA678 : full_adder port map (N2_14_62,N2_15_62,N2_17_62,N3_22_62,N3_23_63);
-- In matrix 2 adding FA to column 63 
	-- signal N3_0_63 : std_logic;
	-- signal N3_1_64 : std_logic;
	FA679 : full_adder port map (N0_32_63,N0_33_63,N0_34_63,N3_0_63,N3_1_64);
-- In matrix 2 adding FA to column 63 
	-- signal N3_2_63 : std_logic;
	-- signal N3_3_64 : std_logic;
	FA680 : full_adder port map (N0_35_63,N0_36_63,N0_37_63,N3_2_63,N3_3_64);
-- In matrix 2 adding FA to column 63 
	-- signal N3_4_63 : std_logic;
	-- signal N3_5_64 : std_logic;
	FA681 : full_adder port map (N0_38_63,N0_39_63,N0_40_63,N3_4_63,N3_5_64);
-- In matrix 2 adding FA to column 63 
	-- signal N3_6_63 : std_logic;
	-- signal N3_7_64 : std_logic;
	FA682 : full_adder port map (N0_41_63,N0_42_63,N0_43_63,N3_6_63,N3_7_64);
-- In matrix 2 adding FA to column 63 
	-- signal N3_8_63 : std_logic;
	-- signal N3_9_64 : std_logic;
	FA683 : full_adder port map (N0_44_63,N0_45_63,N0_46_63,N3_8_63,N3_9_64);
-- In matrix 2 adding FA to column 63 
	-- signal N3_10_63 : std_logic;
	-- signal N3_11_64 : std_logic;
	FA684 : full_adder port map (N0_47_63,N0_48_63,N0_49_63,N3_10_63,N3_11_64);
-- In matrix 2 adding FA to column 63 
	-- signal N3_12_63 : std_logic;
	-- signal N3_13_64 : std_logic;
	FA685 : full_adder port map (N0_50_63,N0_51_63,N0_52_63,N3_12_63,N3_13_64);
-- In matrix 2 adding FA to column 63 
	-- signal N3_14_63 : std_logic;
	-- signal N3_15_64 : std_logic;
	FA686 : full_adder port map (N2_0_63,N2_1_63,N2_2_63,N3_14_63,N3_15_64);
-- In matrix 2 adding FA to column 63 
	-- signal N3_16_63 : std_logic;
	-- signal N3_17_64 : std_logic;
	FA687 : full_adder port map (N2_3_63,N2_4_63,N2_5_63,N3_16_63,N3_17_64);
-- In matrix 2 adding FA to column 63 
	-- signal N3_18_63 : std_logic;
	-- signal N3_19_64 : std_logic;
	FA688 : full_adder port map (N2_6_63,N2_7_63,N2_8_63,N3_18_63,N3_19_64);
-- In matrix 2 adding FA to column 63 
	-- signal N3_20_63 : std_logic;
	-- signal N3_21_64 : std_logic;
	FA689 : full_adder port map (N2_9_63,N2_10_63,N2_11_63,N3_20_63,N3_21_64);
-- In matrix 2 adding FA to column 63 
	-- signal N3_22_63 : std_logic;
	-- signal N3_23_64 : std_logic;
	FA690 : full_adder port map (N2_12_63,N2_13_63,N2_15_63,N3_22_63,N3_23_64);
-- In matrix 2 adding FA to column 64 
	-- signal N3_0_64 : std_logic;
	-- signal N3_1_65 : std_logic;
	FA691 : full_adder port map (N0_30_64,N0_31_64,N0_32_64,N3_0_64,N3_1_65);
-- In matrix 2 adding FA to column 64 
	-- signal N3_2_64 : std_logic;
	-- signal N3_3_65 : std_logic;
	FA692 : full_adder port map (N0_33_64,N0_34_64,N0_35_64,N3_2_64,N3_3_65);
-- In matrix 2 adding FA to column 64 
	-- signal N3_4_64 : std_logic;
	-- signal N3_5_65 : std_logic;
	FA693 : full_adder port map (N0_36_64,N0_37_64,N0_38_64,N3_4_64,N3_5_65);
-- In matrix 2 adding FA to column 64 
	-- signal N3_6_64 : std_logic;
	-- signal N3_7_65 : std_logic;
	FA694 : full_adder port map (N0_39_64,N0_40_64,N0_41_64,N3_6_64,N3_7_65);
-- In matrix 2 adding FA to column 64 
	-- signal N3_8_64 : std_logic;
	-- signal N3_9_65 : std_logic;
	FA695 : full_adder port map (N0_42_64,N0_43_64,N0_44_64,N3_8_64,N3_9_65);
-- In matrix 2 adding FA to column 64 
	-- signal N3_10_64 : std_logic;
	-- signal N3_11_65 : std_logic;
	FA696 : full_adder port map (N0_45_64,N0_46_64,N0_47_64,N3_10_64,N3_11_65);
-- In matrix 2 adding FA to column 64 
	-- signal N3_12_64 : std_logic;
	-- signal N3_13_65 : std_logic;
	FA697 : full_adder port map (N0_48_64,N0_49_64,N0_50_64,N3_12_64,N3_13_65);
-- In matrix 2 adding FA to column 64 
	-- signal N3_14_64 : std_logic;
	-- signal N3_15_65 : std_logic;
	FA698 : full_adder port map (N0_51_64,N0_52_64,N2_0_64,N3_14_64,N3_15_65);
-- In matrix 2 adding FA to column 64 
	-- signal N3_16_64 : std_logic;
	-- signal N3_17_65 : std_logic;
	FA699 : full_adder port map (N2_1_64,N2_2_64,N2_3_64,N3_16_64,N3_17_65);
-- In matrix 2 adding FA to column 64 
	-- signal N3_18_64 : std_logic;
	-- signal N3_19_65 : std_logic;
	FA700 : full_adder port map (N2_4_64,N2_5_64,N2_6_64,N3_18_64,N3_19_65);
-- In matrix 2 adding FA to column 64 
	-- signal N3_20_64 : std_logic;
	-- signal N3_21_65 : std_logic;
	FA701 : full_adder port map (N2_7_64,N2_8_64,N2_9_64,N3_20_64,N3_21_65);
-- In matrix 2 adding FA to column 64 
	-- signal N3_22_64 : std_logic;
	-- signal N3_23_65 : std_logic;
	FA702 : full_adder port map (N2_10_64,N2_11_64,N2_13_64,N3_22_64,N3_23_65);
-- In matrix 2 adding FA to column 65 
	-- signal N3_0_65 : std_logic;
	-- signal N3_1_66 : std_logic;
	FA703 : full_adder port map (N0_28_65,N0_29_65,N0_30_65,N3_0_65,N3_1_66);
-- In matrix 2 adding FA to column 65 
	-- signal N3_2_65 : std_logic;
	-- signal N3_3_66 : std_logic;
	FA704 : full_adder port map (N0_31_65,N0_32_65,N0_33_65,N3_2_65,N3_3_66);
-- In matrix 2 adding FA to column 65 
	-- signal N3_4_65 : std_logic;
	-- signal N3_5_66 : std_logic;
	FA705 : full_adder port map (N0_34_65,N0_35_65,N0_36_65,N3_4_65,N3_5_66);
-- In matrix 2 adding FA to column 65 
	-- signal N3_6_65 : std_logic;
	-- signal N3_7_66 : std_logic;
	FA706 : full_adder port map (N0_37_65,N0_38_65,N0_39_65,N3_6_65,N3_7_66);
-- In matrix 2 adding FA to column 65 
	-- signal N3_8_65 : std_logic;
	-- signal N3_9_66 : std_logic;
	FA707 : full_adder port map (N0_40_65,N0_41_65,N0_42_65,N3_8_65,N3_9_66);
-- In matrix 2 adding FA to column 65 
	-- signal N3_10_65 : std_logic;
	-- signal N3_11_66 : std_logic;
	FA708 : full_adder port map (N0_43_65,N0_44_65,N0_45_65,N3_10_65,N3_11_66);
-- In matrix 2 adding FA to column 65 
	-- signal N3_12_65 : std_logic;
	-- signal N3_13_66 : std_logic;
	FA709 : full_adder port map (N0_46_65,N0_47_65,N0_48_65,N3_12_65,N3_13_66);
-- In matrix 2 adding FA to column 65 
	-- signal N3_14_65 : std_logic;
	-- signal N3_15_66 : std_logic;
	FA710 : full_adder port map (N0_49_65,N0_50_65,N0_51_65,N3_14_65,N3_15_66);
-- In matrix 2 adding FA to column 65 
	-- signal N3_16_65 : std_logic;
	-- signal N3_17_66 : std_logic;
	FA711 : full_adder port map (N0_52_65,N2_0_65,N2_1_65,N3_16_65,N3_17_66);
-- In matrix 2 adding FA to column 65 
	-- signal N3_18_65 : std_logic;
	-- signal N3_19_66 : std_logic;
	FA712 : full_adder port map (N2_2_65,N2_3_65,N2_4_65,N3_18_65,N3_19_66);
-- In matrix 2 adding FA to column 65 
	-- signal N3_20_65 : std_logic;
	-- signal N3_21_66 : std_logic;
	FA713 : full_adder port map (N2_5_65,N2_6_65,N2_7_65,N3_20_65,N3_21_66);
-- In matrix 2 adding FA to column 65 
	-- signal N3_22_65 : std_logic;
	-- signal N3_23_66 : std_logic;
	FA714 : full_adder port map (N2_8_65,N2_9_65,N2_11_65,N3_22_65,N3_23_66);
-- In matrix 2 adding FA to column 66 
	-- signal N3_0_66 : std_logic;
	-- signal N3_1_67 : std_logic;
	FA715 : full_adder port map (N0_26_66,N0_27_66,N0_28_66,N3_0_66,N3_1_67);
-- In matrix 2 adding FA to column 66 
	-- signal N3_2_66 : std_logic;
	-- signal N3_3_67 : std_logic;
	FA716 : full_adder port map (N0_29_66,N0_30_66,N0_31_66,N3_2_66,N3_3_67);
-- In matrix 2 adding FA to column 66 
	-- signal N3_4_66 : std_logic;
	-- signal N3_5_67 : std_logic;
	FA717 : full_adder port map (N0_32_66,N0_33_66,N0_34_66,N3_4_66,N3_5_67);
-- In matrix 2 adding FA to column 66 
	-- signal N3_6_66 : std_logic;
	-- signal N3_7_67 : std_logic;
	FA718 : full_adder port map (N0_35_66,N0_36_66,N0_37_66,N3_6_66,N3_7_67);
-- In matrix 2 adding FA to column 66 
	-- signal N3_8_66 : std_logic;
	-- signal N3_9_67 : std_logic;
	FA719 : full_adder port map (N0_38_66,N0_39_66,N0_40_66,N3_8_66,N3_9_67);
-- In matrix 2 adding FA to column 66 
	-- signal N3_10_66 : std_logic;
	-- signal N3_11_67 : std_logic;
	FA720 : full_adder port map (N0_41_66,N0_42_66,N0_43_66,N3_10_66,N3_11_67);
-- In matrix 2 adding FA to column 66 
	-- signal N3_12_66 : std_logic;
	-- signal N3_13_67 : std_logic;
	FA721 : full_adder port map (N0_44_66,N0_45_66,N0_46_66,N3_12_66,N3_13_67);
-- In matrix 2 adding FA to column 66 
	-- signal N3_14_66 : std_logic;
	-- signal N3_15_67 : std_logic;
	FA722 : full_adder port map (N0_47_66,N0_48_66,N0_49_66,N3_14_66,N3_15_67);
-- In matrix 2 adding FA to column 66 
	-- signal N3_16_66 : std_logic;
	-- signal N3_17_67 : std_logic;
	FA723 : full_adder port map (N0_50_66,N0_51_66,N0_52_66,N3_16_66,N3_17_67);
-- In matrix 2 adding FA to column 66 
	-- signal N3_18_66 : std_logic;
	-- signal N3_19_67 : std_logic;
	FA724 : full_adder port map (N2_0_66,N2_1_66,N2_2_66,N3_18_66,N3_19_67);
-- In matrix 2 adding FA to column 66 
	-- signal N3_20_66 : std_logic;
	-- signal N3_21_67 : std_logic;
	FA725 : full_adder port map (N2_3_66,N2_4_66,N2_5_66,N3_20_66,N3_21_67);
-- In matrix 2 adding FA to column 66 
	-- signal N3_22_66 : std_logic;
	-- signal N3_23_67 : std_logic;
	FA726 : full_adder port map (N2_6_66,N2_7_66,N2_9_66,N3_22_66,N3_23_67);
-- In matrix 2 adding FA to column 67 
	-- signal N3_0_67 : std_logic;
	-- signal N3_1_68 : std_logic;
	FA727 : full_adder port map (N0_24_67,N0_25_67,N0_26_67,N3_0_67,N3_1_68);
-- In matrix 2 adding FA to column 67 
	-- signal N3_2_67 : std_logic;
	-- signal N3_3_68 : std_logic;
	FA728 : full_adder port map (N0_27_67,N0_28_67,N0_29_67,N3_2_67,N3_3_68);
-- In matrix 2 adding FA to column 67 
	-- signal N3_4_67 : std_logic;
	-- signal N3_5_68 : std_logic;
	FA729 : full_adder port map (N0_30_67,N0_31_67,N0_32_67,N3_4_67,N3_5_68);
-- In matrix 2 adding FA to column 67 
	-- signal N3_6_67 : std_logic;
	-- signal N3_7_68 : std_logic;
	FA730 : full_adder port map (N0_33_67,N0_34_67,N0_35_67,N3_6_67,N3_7_68);
-- In matrix 2 adding FA to column 67 
	-- signal N3_8_67 : std_logic;
	-- signal N3_9_68 : std_logic;
	FA731 : full_adder port map (N0_36_67,N0_37_67,N0_38_67,N3_8_67,N3_9_68);
-- In matrix 2 adding FA to column 67 
	-- signal N3_10_67 : std_logic;
	-- signal N3_11_68 : std_logic;
	FA732 : full_adder port map (N0_39_67,N0_40_67,N0_41_67,N3_10_67,N3_11_68);
-- In matrix 2 adding FA to column 67 
	-- signal N3_12_67 : std_logic;
	-- signal N3_13_68 : std_logic;
	FA733 : full_adder port map (N0_42_67,N0_43_67,N0_44_67,N3_12_67,N3_13_68);
-- In matrix 2 adding FA to column 67 
	-- signal N3_14_67 : std_logic;
	-- signal N3_15_68 : std_logic;
	FA734 : full_adder port map (N0_45_67,N0_46_67,N0_47_67,N3_14_67,N3_15_68);
-- In matrix 2 adding FA to column 67 
	-- signal N3_16_67 : std_logic;
	-- signal N3_17_68 : std_logic;
	FA735 : full_adder port map (N0_48_67,N0_49_67,N0_50_67,N3_16_67,N3_17_68);
-- In matrix 2 adding FA to column 67 
	-- signal N3_18_67 : std_logic;
	-- signal N3_19_68 : std_logic;
	FA736 : full_adder port map (N0_51_67,N0_52_67,N2_0_67,N3_18_67,N3_19_68);
-- In matrix 2 adding FA to column 67 
	-- signal N3_20_67 : std_logic;
	-- signal N3_21_68 : std_logic;
	FA737 : full_adder port map (N2_1_67,N2_2_67,N2_3_67,N3_20_67,N3_21_68);
-- In matrix 2 adding FA to column 67 
	-- signal N3_22_67 : std_logic;
	-- signal N3_23_68 : std_logic;
	FA738 : full_adder port map (N2_4_67,N2_5_67,N2_7_67,N3_22_67,N3_23_68);
-- In matrix 2 adding FA to column 68 
	-- signal N3_0_68 : std_logic;
	-- signal N3_1_69 : std_logic;
	FA739 : full_adder port map (N0_22_68,N0_23_68,N0_24_68,N3_0_68,N3_1_69);
-- In matrix 2 adding FA to column 68 
	-- signal N3_2_68 : std_logic;
	-- signal N3_3_69 : std_logic;
	FA740 : full_adder port map (N0_25_68,N0_26_68,N0_27_68,N3_2_68,N3_3_69);
-- In matrix 2 adding FA to column 68 
	-- signal N3_4_68 : std_logic;
	-- signal N3_5_69 : std_logic;
	FA741 : full_adder port map (N0_28_68,N0_29_68,N0_30_68,N3_4_68,N3_5_69);
-- In matrix 2 adding FA to column 68 
	-- signal N3_6_68 : std_logic;
	-- signal N3_7_69 : std_logic;
	FA742 : full_adder port map (N0_31_68,N0_32_68,N0_33_68,N3_6_68,N3_7_69);
-- In matrix 2 adding FA to column 68 
	-- signal N3_8_68 : std_logic;
	-- signal N3_9_69 : std_logic;
	FA743 : full_adder port map (N0_34_68,N0_35_68,N0_36_68,N3_8_68,N3_9_69);
-- In matrix 2 adding FA to column 68 
	-- signal N3_10_68 : std_logic;
	-- signal N3_11_69 : std_logic;
	FA744 : full_adder port map (N0_37_68,N0_38_68,N0_39_68,N3_10_68,N3_11_69);
-- In matrix 2 adding FA to column 68 
	-- signal N3_12_68 : std_logic;
	-- signal N3_13_69 : std_logic;
	FA745 : full_adder port map (N0_40_68,N0_41_68,N0_42_68,N3_12_68,N3_13_69);
-- In matrix 2 adding FA to column 68 
	-- signal N3_14_68 : std_logic;
	-- signal N3_15_69 : std_logic;
	FA746 : full_adder port map (N0_43_68,N0_44_68,N0_45_68,N3_14_68,N3_15_69);
-- In matrix 2 adding FA to column 68 
	-- signal N3_16_68 : std_logic;
	-- signal N3_17_69 : std_logic;
	FA747 : full_adder port map (N0_46_68,N0_47_68,N0_48_68,N3_16_68,N3_17_69);
-- In matrix 2 adding FA to column 68 
	-- signal N3_18_68 : std_logic;
	-- signal N3_19_69 : std_logic;
	FA748 : full_adder port map (N0_49_68,N0_50_68,N0_51_68,N3_18_68,N3_19_69);
-- In matrix 2 adding FA to column 68 
	-- signal N3_20_68 : std_logic;
	-- signal N3_21_69 : std_logic;
	FA749 : full_adder port map (N0_52_68,N2_0_68,N2_1_68,N3_20_68,N3_21_69);
-- In matrix 2 adding FA to column 68 
	-- signal N3_22_68 : std_logic;
	-- signal N3_23_69 : std_logic;
	FA750 : full_adder port map (N2_2_68,N2_3_68,N2_5_68,N3_22_68,N3_23_69);
-- In matrix 2 adding FA to column 69 
	-- signal N3_0_69 : std_logic;
	-- signal N3_1_70 : std_logic;
	FA751 : full_adder port map (N0_20_69,N0_21_69,N0_22_69,N3_0_69,N3_1_70);
-- In matrix 2 adding FA to column 69 
	-- signal N3_2_69 : std_logic;
	-- signal N3_3_70 : std_logic;
	FA752 : full_adder port map (N0_23_69,N0_24_69,N0_25_69,N3_2_69,N3_3_70);
-- In matrix 2 adding FA to column 69 
	-- signal N3_4_69 : std_logic;
	-- signal N3_5_70 : std_logic;
	FA753 : full_adder port map (N0_26_69,N0_27_69,N0_28_69,N3_4_69,N3_5_70);
-- In matrix 2 adding FA to column 69 
	-- signal N3_6_69 : std_logic;
	-- signal N3_7_70 : std_logic;
	FA754 : full_adder port map (N0_29_69,N0_30_69,N0_31_69,N3_6_69,N3_7_70);
-- In matrix 2 adding FA to column 69 
	-- signal N3_8_69 : std_logic;
	-- signal N3_9_70 : std_logic;
	FA755 : full_adder port map (N0_32_69,N0_33_69,N0_34_69,N3_8_69,N3_9_70);
-- In matrix 2 adding FA to column 69 
	-- signal N3_10_69 : std_logic;
	-- signal N3_11_70 : std_logic;
	FA756 : full_adder port map (N0_35_69,N0_36_69,N0_37_69,N3_10_69,N3_11_70);
-- In matrix 2 adding FA to column 69 
	-- signal N3_12_69 : std_logic;
	-- signal N3_13_70 : std_logic;
	FA757 : full_adder port map (N0_38_69,N0_39_69,N0_40_69,N3_12_69,N3_13_70);
-- In matrix 2 adding FA to column 69 
	-- signal N3_14_69 : std_logic;
	-- signal N3_15_70 : std_logic;
	FA758 : full_adder port map (N0_41_69,N0_42_69,N0_43_69,N3_14_69,N3_15_70);
-- In matrix 2 adding FA to column 69 
	-- signal N3_16_69 : std_logic;
	-- signal N3_17_70 : std_logic;
	FA759 : full_adder port map (N0_44_69,N0_45_69,N0_46_69,N3_16_69,N3_17_70);
-- In matrix 2 adding FA to column 69 
	-- signal N3_18_69 : std_logic;
	-- signal N3_19_70 : std_logic;
	FA760 : full_adder port map (N0_47_69,N0_48_69,N0_49_69,N3_18_69,N3_19_70);
-- In matrix 2 adding FA to column 69 
	-- signal N3_20_69 : std_logic;
	-- signal N3_21_70 : std_logic;
	FA761 : full_adder port map (N0_50_69,N0_51_69,N0_52_69,N3_20_69,N3_21_70);
-- In matrix 2 adding FA to column 69 
	-- signal N3_22_69 : std_logic;
	-- signal N3_23_70 : std_logic;
	FA762 : full_adder port map (N2_0_69,N2_1_69,N2_3_69,N3_22_69,N3_23_70);
-- In matrix 2 adding FA to column 70 
	-- signal N3_0_70 : std_logic;
	-- signal N3_1_71 : std_logic;
	FA763 : full_adder port map (N0_18_70,N0_19_70,N0_20_70,N3_0_70,N3_1_71);
-- In matrix 2 adding FA to column 70 
	-- signal N3_2_70 : std_logic;
	-- signal N3_3_71 : std_logic;
	FA764 : full_adder port map (N0_21_70,N0_22_70,N0_23_70,N3_2_70,N3_3_71);
-- In matrix 2 adding FA to column 70 
	-- signal N3_4_70 : std_logic;
	-- signal N3_5_71 : std_logic;
	FA765 : full_adder port map (N0_24_70,N0_25_70,N0_26_70,N3_4_70,N3_5_71);
-- In matrix 2 adding FA to column 70 
	-- signal N3_6_70 : std_logic;
	-- signal N3_7_71 : std_logic;
	FA766 : full_adder port map (N0_27_70,N0_28_70,N0_29_70,N3_6_70,N3_7_71);
-- In matrix 2 adding FA to column 70 
	-- signal N3_8_70 : std_logic;
	-- signal N3_9_71 : std_logic;
	FA767 : full_adder port map (N0_30_70,N0_31_70,N0_32_70,N3_8_70,N3_9_71);
-- In matrix 2 adding FA to column 70 
	-- signal N3_10_70 : std_logic;
	-- signal N3_11_71 : std_logic;
	FA768 : full_adder port map (N0_33_70,N0_34_70,N0_35_70,N3_10_70,N3_11_71);
-- In matrix 2 adding FA to column 70 
	-- signal N3_12_70 : std_logic;
	-- signal N3_13_71 : std_logic;
	FA769 : full_adder port map (N0_36_70,N0_37_70,N0_38_70,N3_12_70,N3_13_71);
-- In matrix 2 adding FA to column 70 
	-- signal N3_14_70 : std_logic;
	-- signal N3_15_71 : std_logic;
	FA770 : full_adder port map (N0_39_70,N0_40_70,N0_41_70,N3_14_70,N3_15_71);
-- In matrix 2 adding FA to column 70 
	-- signal N3_16_70 : std_logic;
	-- signal N3_17_71 : std_logic;
	FA771 : full_adder port map (N0_42_70,N0_43_70,N0_44_70,N3_16_70,N3_17_71);
-- In matrix 2 adding FA to column 70 
	-- signal N3_18_70 : std_logic;
	-- signal N3_19_71 : std_logic;
	FA772 : full_adder port map (N0_45_70,N0_46_70,N0_47_70,N3_18_70,N3_19_71);
-- In matrix 2 adding FA to column 70 
	-- signal N3_20_70 : std_logic;
	-- signal N3_21_71 : std_logic;
	FA773 : full_adder port map (N0_48_70,N0_49_70,N0_50_70,N3_20_70,N3_21_71);
-- In matrix 2 adding FA to column 70 
	-- signal N3_22_70 : std_logic;
	-- signal N3_23_71 : std_logic;
	FA774 : full_adder port map (N0_51_70,N0_52_70,N2_1_70,N3_22_70,N3_23_71);
-- In matrix 2 adding FA to column 71 
	-- signal N3_0_71 : std_logic;
	-- signal N3_1_72 : std_logic;
	FA775 : full_adder port map (N0_19_71,N0_20_71,N0_21_71,N3_0_71,N3_1_72);
-- In matrix 2 adding FA to column 71 
	-- signal N3_2_71 : std_logic;
	-- signal N3_3_72 : std_logic;
	FA776 : full_adder port map (N0_22_71,N0_23_71,N0_24_71,N3_2_71,N3_3_72);
-- In matrix 2 adding FA to column 71 
	-- signal N3_4_71 : std_logic;
	-- signal N3_5_72 : std_logic;
	FA777 : full_adder port map (N0_25_71,N0_26_71,N0_27_71,N3_4_71,N3_5_72);
-- In matrix 2 adding FA to column 71 
	-- signal N3_6_71 : std_logic;
	-- signal N3_7_72 : std_logic;
	FA778 : full_adder port map (N0_28_71,N0_29_71,N0_30_71,N3_6_71,N3_7_72);
-- In matrix 2 adding FA to column 71 
	-- signal N3_8_71 : std_logic;
	-- signal N3_9_72 : std_logic;
	FA779 : full_adder port map (N0_31_71,N0_32_71,N0_33_71,N3_8_71,N3_9_72);
-- In matrix 2 adding FA to column 71 
	-- signal N3_10_71 : std_logic;
	-- signal N3_11_72 : std_logic;
	FA780 : full_adder port map (N0_34_71,N0_35_71,N0_36_71,N3_10_71,N3_11_72);
-- In matrix 2 adding FA to column 71 
	-- signal N3_12_71 : std_logic;
	-- signal N3_13_72 : std_logic;
	FA781 : full_adder port map (N0_37_71,N0_38_71,N0_39_71,N3_12_71,N3_13_72);
-- In matrix 2 adding FA to column 71 
	-- signal N3_14_71 : std_logic;
	-- signal N3_15_72 : std_logic;
	FA782 : full_adder port map (N0_40_71,N0_41_71,N0_42_71,N3_14_71,N3_15_72);
-- In matrix 2 adding FA to column 71 
	-- signal N3_16_71 : std_logic;
	-- signal N3_17_72 : std_logic;
	FA783 : full_adder port map (N0_43_71,N0_44_71,N0_45_71,N3_16_71,N3_17_72);
-- In matrix 2 adding FA to column 71 
	-- signal N3_18_71 : std_logic;
	-- signal N3_19_72 : std_logic;
	FA784 : full_adder port map (N0_46_71,N0_47_71,N0_48_71,N3_18_71,N3_19_72);
-- In matrix 2 adding FA to column 71 
	-- signal N3_20_71 : std_logic;
	-- signal N3_21_72 : std_logic;
	FA785 : full_adder port map (N0_49_71,N0_50_71,N0_51_71,N3_20_71,N3_21_72);
-- In matrix 2 adding FA to column 72 
	-- signal N3_0_72 : std_logic;
	-- signal N3_1_73 : std_logic;
	FA786 : full_adder port map (N0_20_72,N0_21_72,N0_22_72,N3_0_72,N3_1_73);
-- In matrix 2 adding FA to column 72 
	-- signal N3_2_72 : std_logic;
	-- signal N3_3_73 : std_logic;
	FA787 : full_adder port map (N0_23_72,N0_24_72,N0_25_72,N3_2_72,N3_3_73);
-- In matrix 2 adding FA to column 72 
	-- signal N3_4_72 : std_logic;
	-- signal N3_5_73 : std_logic;
	FA788 : full_adder port map (N0_26_72,N0_27_72,N0_28_72,N3_4_72,N3_5_73);
-- In matrix 2 adding FA to column 72 
	-- signal N3_6_72 : std_logic;
	-- signal N3_7_73 : std_logic;
	FA789 : full_adder port map (N0_29_72,N0_30_72,N0_31_72,N3_6_72,N3_7_73);
-- In matrix 2 adding FA to column 72 
	-- signal N3_8_72 : std_logic;
	-- signal N3_9_73 : std_logic;
	FA790 : full_adder port map (N0_32_72,N0_33_72,N0_34_72,N3_8_72,N3_9_73);
-- In matrix 2 adding FA to column 72 
	-- signal N3_10_72 : std_logic;
	-- signal N3_11_73 : std_logic;
	FA791 : full_adder port map (N0_35_72,N0_36_72,N0_37_72,N3_10_72,N3_11_73);
-- In matrix 2 adding FA to column 72 
	-- signal N3_12_72 : std_logic;
	-- signal N3_13_73 : std_logic;
	FA792 : full_adder port map (N0_38_72,N0_39_72,N0_40_72,N3_12_72,N3_13_73);
-- In matrix 2 adding FA to column 72 
	-- signal N3_14_72 : std_logic;
	-- signal N3_15_73 : std_logic;
	FA793 : full_adder port map (N0_41_72,N0_42_72,N0_43_72,N3_14_72,N3_15_73);
-- In matrix 2 adding FA to column 72 
	-- signal N3_16_72 : std_logic;
	-- signal N3_17_73 : std_logic;
	FA794 : full_adder port map (N0_44_72,N0_45_72,N0_46_72,N3_16_72,N3_17_73);
-- In matrix 2 adding FA to column 72 
	-- signal N3_18_72 : std_logic;
	-- signal N3_19_73 : std_logic;
	FA795 : full_adder port map (N0_47_72,N0_48_72,N0_49_72,N3_18_72,N3_19_73);
-- In matrix 2 adding FA to column 73 
	-- signal N3_0_73 : std_logic;
	-- signal N3_1_74 : std_logic;
	FA796 : full_adder port map (N0_21_73,N0_22_73,N0_23_73,N3_0_73,N3_1_74);
-- In matrix 2 adding FA to column 73 
	-- signal N3_2_73 : std_logic;
	-- signal N3_3_74 : std_logic;
	FA797 : full_adder port map (N0_24_73,N0_25_73,N0_26_73,N3_2_73,N3_3_74);
-- In matrix 2 adding FA to column 73 
	-- signal N3_4_73 : std_logic;
	-- signal N3_5_74 : std_logic;
	FA798 : full_adder port map (N0_27_73,N0_28_73,N0_29_73,N3_4_73,N3_5_74);
-- In matrix 2 adding FA to column 73 
	-- signal N3_6_73 : std_logic;
	-- signal N3_7_74 : std_logic;
	FA799 : full_adder port map (N0_30_73,N0_31_73,N0_32_73,N3_6_73,N3_7_74);
-- In matrix 2 adding FA to column 73 
	-- signal N3_8_73 : std_logic;
	-- signal N3_9_74 : std_logic;
	FA800 : full_adder port map (N0_33_73,N0_34_73,N0_35_73,N3_8_73,N3_9_74);
-- In matrix 2 adding FA to column 73 
	-- signal N3_10_73 : std_logic;
	-- signal N3_11_74 : std_logic;
	FA801 : full_adder port map (N0_36_73,N0_37_73,N0_38_73,N3_10_73,N3_11_74);
-- In matrix 2 adding FA to column 73 
	-- signal N3_12_73 : std_logic;
	-- signal N3_13_74 : std_logic;
	FA802 : full_adder port map (N0_39_73,N0_40_73,N0_41_73,N3_12_73,N3_13_74);
-- In matrix 2 adding FA to column 73 
	-- signal N3_14_73 : std_logic;
	-- signal N3_15_74 : std_logic;
	FA803 : full_adder port map (N0_42_73,N0_43_73,N0_44_73,N3_14_73,N3_15_74);
-- In matrix 2 adding FA to column 73 
	-- signal N3_16_73 : std_logic;
	-- signal N3_17_74 : std_logic;
	FA804 : full_adder port map (N0_45_73,N0_46_73,N0_47_73,N3_16_73,N3_17_74);
-- In matrix 2 adding FA to column 74 
	-- signal N3_0_74 : std_logic;
	-- signal N3_1_75 : std_logic;
	FA805 : full_adder port map (N0_22_74,N0_23_74,N0_24_74,N3_0_74,N3_1_75);
-- In matrix 2 adding FA to column 74 
	-- signal N3_2_74 : std_logic;
	-- signal N3_3_75 : std_logic;
	FA806 : full_adder port map (N0_25_74,N0_26_74,N0_27_74,N3_2_74,N3_3_75);
-- In matrix 2 adding FA to column 74 
	-- signal N3_4_74 : std_logic;
	-- signal N3_5_75 : std_logic;
	FA807 : full_adder port map (N0_28_74,N0_29_74,N0_30_74,N3_4_74,N3_5_75);
-- In matrix 2 adding FA to column 74 
	-- signal N3_6_74 : std_logic;
	-- signal N3_7_75 : std_logic;
	FA808 : full_adder port map (N0_31_74,N0_32_74,N0_33_74,N3_6_74,N3_7_75);
-- In matrix 2 adding FA to column 74 
	-- signal N3_8_74 : std_logic;
	-- signal N3_9_75 : std_logic;
	FA809 : full_adder port map (N0_34_74,N0_35_74,N0_36_74,N3_8_74,N3_9_75);
-- In matrix 2 adding FA to column 74 
	-- signal N3_10_74 : std_logic;
	-- signal N3_11_75 : std_logic;
	FA810 : full_adder port map (N0_37_74,N0_38_74,N0_39_74,N3_10_74,N3_11_75);
-- In matrix 2 adding FA to column 74 
	-- signal N3_12_74 : std_logic;
	-- signal N3_13_75 : std_logic;
	FA811 : full_adder port map (N0_40_74,N0_41_74,N0_42_74,N3_12_74,N3_13_75);
-- In matrix 2 adding FA to column 74 
	-- signal N3_14_74 : std_logic;
	-- signal N3_15_75 : std_logic;
	FA812 : full_adder port map (N0_43_74,N0_44_74,N0_45_74,N3_14_74,N3_15_75);
-- In matrix 2 adding FA to column 75 
	-- signal N3_0_75 : std_logic;
	-- signal N3_1_76 : std_logic;
	FA813 : full_adder port map (N0_23_75,N0_24_75,N0_25_75,N3_0_75,N3_1_76);
-- In matrix 2 adding FA to column 75 
	-- signal N3_2_75 : std_logic;
	-- signal N3_3_76 : std_logic;
	FA814 : full_adder port map (N0_26_75,N0_27_75,N0_28_75,N3_2_75,N3_3_76);
-- In matrix 2 adding FA to column 75 
	-- signal N3_4_75 : std_logic;
	-- signal N3_5_76 : std_logic;
	FA815 : full_adder port map (N0_29_75,N0_30_75,N0_31_75,N3_4_75,N3_5_76);
-- In matrix 2 adding FA to column 75 
	-- signal N3_6_75 : std_logic;
	-- signal N3_7_76 : std_logic;
	FA816 : full_adder port map (N0_32_75,N0_33_75,N0_34_75,N3_6_75,N3_7_76);
-- In matrix 2 adding FA to column 75 
	-- signal N3_8_75 : std_logic;
	-- signal N3_9_76 : std_logic;
	FA817 : full_adder port map (N0_35_75,N0_36_75,N0_37_75,N3_8_75,N3_9_76);
-- In matrix 2 adding FA to column 75 
	-- signal N3_10_75 : std_logic;
	-- signal N3_11_76 : std_logic;
	FA818 : full_adder port map (N0_38_75,N0_39_75,N0_40_75,N3_10_75,N3_11_76);
-- In matrix 2 adding FA to column 75 
	-- signal N3_12_75 : std_logic;
	-- signal N3_13_76 : std_logic;
	FA819 : full_adder port map (N0_41_75,N0_42_75,N0_43_75,N3_12_75,N3_13_76);
-- In matrix 2 adding FA to column 76 
	-- signal N3_0_76 : std_logic;
	-- signal N3_1_77 : std_logic;
	FA820 : full_adder port map (N0_24_76,N0_25_76,N0_26_76,N3_0_76,N3_1_77);
-- In matrix 2 adding FA to column 76 
	-- signal N3_2_76 : std_logic;
	-- signal N3_3_77 : std_logic;
	FA821 : full_adder port map (N0_27_76,N0_28_76,N0_29_76,N3_2_76,N3_3_77);
-- In matrix 2 adding FA to column 76 
	-- signal N3_4_76 : std_logic;
	-- signal N3_5_77 : std_logic;
	FA822 : full_adder port map (N0_30_76,N0_31_76,N0_32_76,N3_4_76,N3_5_77);
-- In matrix 2 adding FA to column 76 
	-- signal N3_6_76 : std_logic;
	-- signal N3_7_77 : std_logic;
	FA823 : full_adder port map (N0_33_76,N0_34_76,N0_35_76,N3_6_76,N3_7_77);
-- In matrix 2 adding FA to column 76 
	-- signal N3_8_76 : std_logic;
	-- signal N3_9_77 : std_logic;
	FA824 : full_adder port map (N0_36_76,N0_37_76,N0_38_76,N3_8_76,N3_9_77);
-- In matrix 2 adding FA to column 76 
	-- signal N3_10_76 : std_logic;
	-- signal N3_11_77 : std_logic;
	FA825 : full_adder port map (N0_39_76,N0_40_76,N0_41_76,N3_10_76,N3_11_77);
-- In matrix 2 adding FA to column 77 
	-- signal N3_0_77 : std_logic;
	-- signal N3_1_78 : std_logic;
	FA826 : full_adder port map (N0_25_77,N0_26_77,N0_27_77,N3_0_77,N3_1_78);
-- In matrix 2 adding FA to column 77 
	-- signal N3_2_77 : std_logic;
	-- signal N3_3_78 : std_logic;
	FA827 : full_adder port map (N0_28_77,N0_29_77,N0_30_77,N3_2_77,N3_3_78);
-- In matrix 2 adding FA to column 77 
	-- signal N3_4_77 : std_logic;
	-- signal N3_5_78 : std_logic;
	FA828 : full_adder port map (N0_31_77,N0_32_77,N0_33_77,N3_4_77,N3_5_78);
-- In matrix 2 adding FA to column 77 
	-- signal N3_6_77 : std_logic;
	-- signal N3_7_78 : std_logic;
	FA829 : full_adder port map (N0_34_77,N0_35_77,N0_36_77,N3_6_77,N3_7_78);
-- In matrix 2 adding FA to column 77 
	-- signal N3_8_77 : std_logic;
	-- signal N3_9_78 : std_logic;
	FA830 : full_adder port map (N0_37_77,N0_38_77,N0_39_77,N3_8_77,N3_9_78);
-- In matrix 2 adding FA to column 78 
	-- signal N3_0_78 : std_logic;
	-- signal N3_1_79 : std_logic;
	FA831 : full_adder port map (N0_26_78,N0_27_78,N0_28_78,N3_0_78,N3_1_79);
-- In matrix 2 adding FA to column 78 
	-- signal N3_2_78 : std_logic;
	-- signal N3_3_79 : std_logic;
	FA832 : full_adder port map (N0_29_78,N0_30_78,N0_31_78,N3_2_78,N3_3_79);
-- In matrix 2 adding FA to column 78 
	-- signal N3_4_78 : std_logic;
	-- signal N3_5_79 : std_logic;
	FA833 : full_adder port map (N0_32_78,N0_33_78,N0_34_78,N3_4_78,N3_5_79);
-- In matrix 2 adding FA to column 78 
	-- signal N3_6_78 : std_logic;
	-- signal N3_7_79 : std_logic;
	FA834 : full_adder port map (N0_35_78,N0_36_78,N0_37_78,N3_6_78,N3_7_79);
-- In matrix 2 adding FA to column 79 
	-- signal N3_0_79 : std_logic;
	-- signal N3_1_80 : std_logic;
	FA835 : full_adder port map (N0_27_79,N0_28_79,N0_29_79,N3_0_79,N3_1_80);
-- In matrix 2 adding FA to column 79 
	-- signal N3_2_79 : std_logic;
	-- signal N3_3_80 : std_logic;
	FA836 : full_adder port map (N0_30_79,N0_31_79,N0_32_79,N3_2_79,N3_3_80);
-- In matrix 2 adding FA to column 79 
	-- signal N3_4_79 : std_logic;
	-- signal N3_5_80 : std_logic;
	FA837 : full_adder port map (N0_33_79,N0_34_79,N0_35_79,N3_4_79,N3_5_80);
-- In matrix 2 adding FA to column 80 
	-- signal N3_0_80 : std_logic;
	-- signal N3_1_81 : std_logic;
	FA838 : full_adder port map (N0_28_80,N0_29_80,N0_30_80,N3_0_80,N3_1_81);
-- In matrix 2 adding FA to column 80 
	-- signal N3_2_80 : std_logic;
	-- signal N3_3_81 : std_logic;
	FA839 : full_adder port map (N0_31_80,N0_32_80,N0_33_80,N3_2_80,N3_3_81);
-- In matrix 2 adding FA to column 81 
	-- signal N3_0_81 : std_logic;
	-- signal N3_1_82 : std_logic;
	FA840 : full_adder port map (N0_29_81,N0_30_81,N0_31_81,N3_0_81,N3_1_82);
	-- Elements from matrix 3 
-- In matrix 3 adding HA to column 16 
	-- signal N4_0_16 : std_logic;
	-- signal N4_1_17 : std_logic;
	HA31 : half_adder port map (N0_0_16,N0_1_16,N4_0_16,N4_1_17);
-- In matrix 3 adding FA to column 17 
	-- signal N4_0_17 : std_logic;
	-- signal N4_1_18 : std_logic;
	FA841 : full_adder port map (N0_0_17,N0_1_17,N0_2_17,N4_0_17,N4_1_18);
-- In matrix 3 adding HA to column 17 
	-- signal N4_2_17 : std_logic;
	-- signal N4_3_18 : std_logic;
	HA32 : half_adder port map (N0_3_17,N0_4_17,N4_2_17,N4_3_18);
-- In matrix 3 adding FA to column 18 
	-- signal N4_0_18 : std_logic;
	-- signal N4_1_19 : std_logic;
	FA842 : full_adder port map (N0_0_18,N0_1_18,N0_2_18,N4_0_18,N4_1_19);
-- In matrix 3 adding FA to column 18 
	-- signal N4_2_18 : std_logic;
	-- signal N4_3_19 : std_logic;
	FA843 : full_adder port map (N0_3_18,N0_4_18,N0_5_18,N4_2_18,N4_3_19);
-- In matrix 3 adding HA to column 18 
	-- signal N4_4_18 : std_logic;
	-- signal N4_5_19 : std_logic;
	HA33 : half_adder port map (N0_6_18,N0_7_18,N4_4_18,N4_5_19);
-- In matrix 3 adding FA to column 19 
	-- signal N4_0_19 : std_logic;
	-- signal N4_1_20 : std_logic;
	FA844 : full_adder port map (N0_0_19,N0_1_19,N0_2_19,N4_0_19,N4_1_20);
-- In matrix 3 adding FA to column 19 
	-- signal N4_2_19 : std_logic;
	-- signal N4_3_20 : std_logic;
	FA845 : full_adder port map (N0_3_19,N0_4_19,N0_5_19,N4_2_19,N4_3_20);
-- In matrix 3 adding FA to column 19 
	-- signal N4_4_19 : std_logic;
	-- signal N4_5_20 : std_logic;
	FA846 : full_adder port map (N0_6_19,N0_7_19,N0_8_19,N4_4_19,N4_5_20);
-- In matrix 3 adding HA to column 19 
	-- signal N4_6_19 : std_logic;
	-- signal N4_7_20 : std_logic;
	HA34 : half_adder port map (N0_9_19,N0_10_19,N4_6_19,N4_7_20);
-- In matrix 3 adding FA to column 20 
	-- signal N4_0_20 : std_logic;
	-- signal N4_1_21 : std_logic;
	FA847 : full_adder port map (N0_0_20,N0_1_20,N0_2_20,N4_0_20,N4_1_21);
-- In matrix 3 adding FA to column 20 
	-- signal N4_2_20 : std_logic;
	-- signal N4_3_21 : std_logic;
	FA848 : full_adder port map (N0_3_20,N0_4_20,N0_5_20,N4_2_20,N4_3_21);
-- In matrix 3 adding FA to column 20 
	-- signal N4_4_20 : std_logic;
	-- signal N4_5_21 : std_logic;
	FA849 : full_adder port map (N0_6_20,N0_7_20,N0_8_20,N4_4_20,N4_5_21);
-- In matrix 3 adding FA to column 20 
	-- signal N4_6_20 : std_logic;
	-- signal N4_7_21 : std_logic;
	FA850 : full_adder port map (N0_9_20,N0_10_20,N0_11_20,N4_6_20,N4_7_21);
-- In matrix 3 adding HA to column 20 
	-- signal N4_8_20 : std_logic;
	-- signal N4_9_21 : std_logic;
	HA35 : half_adder port map (N0_12_20,N0_13_20,N4_8_20,N4_9_21);
-- In matrix 3 adding FA to column 21 
	-- signal N4_0_21 : std_logic;
	-- signal N4_1_22 : std_logic;
	FA851 : full_adder port map (N0_0_21,N0_1_21,N0_2_21,N4_0_21,N4_1_22);
-- In matrix 3 adding FA to column 21 
	-- signal N4_2_21 : std_logic;
	-- signal N4_3_22 : std_logic;
	FA852 : full_adder port map (N0_3_21,N0_4_21,N0_5_21,N4_2_21,N4_3_22);
-- In matrix 3 adding FA to column 21 
	-- signal N4_4_21 : std_logic;
	-- signal N4_5_22 : std_logic;
	FA853 : full_adder port map (N0_6_21,N0_7_21,N0_8_21,N4_4_21,N4_5_22);
-- In matrix 3 adding FA to column 21 
	-- signal N4_6_21 : std_logic;
	-- signal N4_7_22 : std_logic;
	FA854 : full_adder port map (N0_9_21,N0_10_21,N0_11_21,N4_6_21,N4_7_22);
-- In matrix 3 adding FA to column 21 
	-- signal N4_8_21 : std_logic;
	-- signal N4_9_22 : std_logic;
	FA855 : full_adder port map (N0_12_21,N0_13_21,N0_14_21,N4_8_21,N4_9_22);
-- In matrix 3 adding HA to column 21 
	-- signal N4_10_21 : std_logic;
	-- signal N4_11_22 : std_logic;
	HA36 : half_adder port map (N0_15_21,N0_16_21,N4_10_21,N4_11_22);
-- In matrix 3 adding FA to column 22 
	-- signal N4_0_22 : std_logic;
	-- signal N4_1_23 : std_logic;
	FA856 : full_adder port map (N0_0_22,N0_1_22,N0_2_22,N4_0_22,N4_1_23);
-- In matrix 3 adding FA to column 22 
	-- signal N4_2_22 : std_logic;
	-- signal N4_3_23 : std_logic;
	FA857 : full_adder port map (N0_3_22,N0_4_22,N0_5_22,N4_2_22,N4_3_23);
-- In matrix 3 adding FA to column 22 
	-- signal N4_4_22 : std_logic;
	-- signal N4_5_23 : std_logic;
	FA858 : full_adder port map (N0_6_22,N0_7_22,N0_8_22,N4_4_22,N4_5_23);
-- In matrix 3 adding FA to column 22 
	-- signal N4_6_22 : std_logic;
	-- signal N4_7_23 : std_logic;
	FA859 : full_adder port map (N0_9_22,N0_10_22,N0_11_22,N4_6_22,N4_7_23);
-- In matrix 3 adding FA to column 22 
	-- signal N4_8_22 : std_logic;
	-- signal N4_9_23 : std_logic;
	FA860 : full_adder port map (N0_12_22,N0_13_22,N0_14_22,N4_8_22,N4_9_23);
-- In matrix 3 adding FA to column 22 
	-- signal N4_10_22 : std_logic;
	-- signal N4_11_23 : std_logic;
	FA861 : full_adder port map (N0_15_22,N0_16_22,N0_17_22,N4_10_22,N4_11_23);
-- In matrix 3 adding HA to column 22 
	-- signal N4_12_22 : std_logic;
	-- signal N4_13_23 : std_logic;
	HA37 : half_adder port map (N0_18_22,N0_19_22,N4_12_22,N4_13_23);
-- In matrix 3 adding FA to column 23 
	-- signal N4_0_23 : std_logic;
	-- signal N4_1_24 : std_logic;
	FA862 : full_adder port map (N0_0_23,N0_1_23,N0_2_23,N4_0_23,N4_1_24);
-- In matrix 3 adding FA to column 23 
	-- signal N4_2_23 : std_logic;
	-- signal N4_3_24 : std_logic;
	FA863 : full_adder port map (N0_3_23,N0_4_23,N0_5_23,N4_2_23,N4_3_24);
-- In matrix 3 adding FA to column 23 
	-- signal N4_4_23 : std_logic;
	-- signal N4_5_24 : std_logic;
	FA864 : full_adder port map (N0_6_23,N0_7_23,N0_8_23,N4_4_23,N4_5_24);
-- In matrix 3 adding FA to column 23 
	-- signal N4_6_23 : std_logic;
	-- signal N4_7_24 : std_logic;
	FA865 : full_adder port map (N0_9_23,N0_10_23,N0_11_23,N4_6_23,N4_7_24);
-- In matrix 3 adding FA to column 23 
	-- signal N4_8_23 : std_logic;
	-- signal N4_9_24 : std_logic;
	FA866 : full_adder port map (N0_12_23,N0_13_23,N0_14_23,N4_8_23,N4_9_24);
-- In matrix 3 adding FA to column 23 
	-- signal N4_10_23 : std_logic;
	-- signal N4_11_24 : std_logic;
	FA867 : full_adder port map (N0_15_23,N0_16_23,N0_17_23,N4_10_23,N4_11_24);
-- In matrix 3 adding FA to column 23 
	-- signal N4_12_23 : std_logic;
	-- signal N4_13_24 : std_logic;
	FA868 : full_adder port map (N0_18_23,N0_19_23,N0_20_23,N4_12_23,N4_13_24);
-- In matrix 3 adding HA to column 23 
	-- signal N4_14_23 : std_logic;
	-- signal N4_15_24 : std_logic;
	HA38 : half_adder port map (N0_21_23,N0_22_23,N4_14_23,N4_15_24);
-- In matrix 3 adding FA to column 24 
	-- signal N4_0_24 : std_logic;
	-- signal N4_1_25 : std_logic;
	FA869 : full_adder port map (N0_2_24,N0_3_24,N0_4_24,N4_0_24,N4_1_25);
-- In matrix 3 adding FA to column 24 
	-- signal N4_2_24 : std_logic;
	-- signal N4_3_25 : std_logic;
	FA870 : full_adder port map (N0_5_24,N0_6_24,N0_7_24,N4_2_24,N4_3_25);
-- In matrix 3 adding FA to column 24 
	-- signal N4_4_24 : std_logic;
	-- signal N4_5_25 : std_logic;
	FA871 : full_adder port map (N0_8_24,N0_9_24,N0_10_24,N4_4_24,N4_5_25);
-- In matrix 3 adding FA to column 24 
	-- signal N4_6_24 : std_logic;
	-- signal N4_7_25 : std_logic;
	FA872 : full_adder port map (N0_11_24,N0_12_24,N0_13_24,N4_6_24,N4_7_25);
-- In matrix 3 adding FA to column 24 
	-- signal N4_8_24 : std_logic;
	-- signal N4_9_25 : std_logic;
	FA873 : full_adder port map (N0_14_24,N0_15_24,N0_16_24,N4_8_24,N4_9_25);
-- In matrix 3 adding FA to column 24 
	-- signal N4_10_24 : std_logic;
	-- signal N4_11_25 : std_logic;
	FA874 : full_adder port map (N0_17_24,N0_18_24,N0_19_24,N4_10_24,N4_11_25);
-- In matrix 3 adding FA to column 24 
	-- signal N4_12_24 : std_logic;
	-- signal N4_13_25 : std_logic;
	FA875 : full_adder port map (N0_20_24,N0_21_24,N0_22_24,N4_12_24,N4_13_25);
-- In matrix 3 adding FA to column 24 
	-- signal N4_14_24 : std_logic;
	-- signal N4_15_25 : std_logic;
	FA876 : full_adder port map (N0_23_24,N0_24_24,N3_0_24,N4_14_24,N4_15_25);
-- In matrix 3 adding FA to column 25 
	-- signal N4_0_25 : std_logic;
	-- signal N4_1_26 : std_logic;
	FA877 : full_adder port map (N0_5_25,N0_6_25,N0_7_25,N4_0_25,N4_1_26);
-- In matrix 3 adding FA to column 25 
	-- signal N4_2_25 : std_logic;
	-- signal N4_3_26 : std_logic;
	FA878 : full_adder port map (N0_8_25,N0_9_25,N0_10_25,N4_2_25,N4_3_26);
-- In matrix 3 adding FA to column 25 
	-- signal N4_4_25 : std_logic;
	-- signal N4_5_26 : std_logic;
	FA879 : full_adder port map (N0_11_25,N0_12_25,N0_13_25,N4_4_25,N4_5_26);
-- In matrix 3 adding FA to column 25 
	-- signal N4_6_25 : std_logic;
	-- signal N4_7_26 : std_logic;
	FA880 : full_adder port map (N0_14_25,N0_15_25,N0_16_25,N4_6_25,N4_7_26);
-- In matrix 3 adding FA to column 25 
	-- signal N4_8_25 : std_logic;
	-- signal N4_9_26 : std_logic;
	FA881 : full_adder port map (N0_17_25,N0_18_25,N0_19_25,N4_8_25,N4_9_26);
-- In matrix 3 adding FA to column 25 
	-- signal N4_10_25 : std_logic;
	-- signal N4_11_26 : std_logic;
	FA882 : full_adder port map (N0_20_25,N0_21_25,N0_22_25,N4_10_25,N4_11_26);
-- In matrix 3 adding FA to column 25 
	-- signal N4_12_25 : std_logic;
	-- signal N4_13_26 : std_logic;
	FA883 : full_adder port map (N0_23_25,N0_24_25,N0_25_25,N4_12_25,N4_13_26);
-- In matrix 3 adding FA to column 25 
	-- signal N4_14_25 : std_logic;
	-- signal N4_15_26 : std_logic;
	FA884 : full_adder port map (N3_0_25,N3_1_25,N3_2_25,N4_14_25,N4_15_26);
-- In matrix 3 adding FA to column 26 
	-- signal N4_0_26 : std_logic;
	-- signal N4_1_27 : std_logic;
	FA885 : full_adder port map (N0_8_26,N0_9_26,N0_10_26,N4_0_26,N4_1_27);
-- In matrix 3 adding FA to column 26 
	-- signal N4_2_26 : std_logic;
	-- signal N4_3_27 : std_logic;
	FA886 : full_adder port map (N0_11_26,N0_12_26,N0_13_26,N4_2_26,N4_3_27);
-- In matrix 3 adding FA to column 26 
	-- signal N4_4_26 : std_logic;
	-- signal N4_5_27 : std_logic;
	FA887 : full_adder port map (N0_14_26,N0_15_26,N0_16_26,N4_4_26,N4_5_27);
-- In matrix 3 adding FA to column 26 
	-- signal N4_6_26 : std_logic;
	-- signal N4_7_27 : std_logic;
	FA888 : full_adder port map (N0_17_26,N0_18_26,N0_19_26,N4_6_26,N4_7_27);
-- In matrix 3 adding FA to column 26 
	-- signal N4_8_26 : std_logic;
	-- signal N4_9_27 : std_logic;
	FA889 : full_adder port map (N0_20_26,N0_21_26,N0_22_26,N4_8_26,N4_9_27);
-- In matrix 3 adding FA to column 26 
	-- signal N4_10_26 : std_logic;
	-- signal N4_11_27 : std_logic;
	FA890 : full_adder port map (N0_23_26,N0_24_26,N0_25_26,N4_10_26,N4_11_27);
-- In matrix 3 adding FA to column 26 
	-- signal N4_12_26 : std_logic;
	-- signal N4_13_27 : std_logic;
	FA891 : full_adder port map (N0_26_26,N3_0_26,N3_1_26,N4_12_26,N4_13_27);
-- In matrix 3 adding FA to column 26 
	-- signal N4_14_26 : std_logic;
	-- signal N4_15_27 : std_logic;
	FA892 : full_adder port map (N3_2_26,N3_3_26,N3_4_26,N4_14_26,N4_15_27);
-- In matrix 3 adding FA to column 27 
	-- signal N4_0_27 : std_logic;
	-- signal N4_1_28 : std_logic;
	FA893 : full_adder port map (N0_11_27,N0_12_27,N0_13_27,N4_0_27,N4_1_28);
-- In matrix 3 adding FA to column 27 
	-- signal N4_2_27 : std_logic;
	-- signal N4_3_28 : std_logic;
	FA894 : full_adder port map (N0_14_27,N0_15_27,N0_16_27,N4_2_27,N4_3_28);
-- In matrix 3 adding FA to column 27 
	-- signal N4_4_27 : std_logic;
	-- signal N4_5_28 : std_logic;
	FA895 : full_adder port map (N0_17_27,N0_18_27,N0_19_27,N4_4_27,N4_5_28);
-- In matrix 3 adding FA to column 27 
	-- signal N4_6_27 : std_logic;
	-- signal N4_7_28 : std_logic;
	FA896 : full_adder port map (N0_20_27,N0_21_27,N0_22_27,N4_6_27,N4_7_28);
-- In matrix 3 adding FA to column 27 
	-- signal N4_8_27 : std_logic;
	-- signal N4_9_28 : std_logic;
	FA897 : full_adder port map (N0_23_27,N0_24_27,N0_25_27,N4_8_27,N4_9_28);
-- In matrix 3 adding FA to column 27 
	-- signal N4_10_27 : std_logic;
	-- signal N4_11_28 : std_logic;
	FA898 : full_adder port map (N0_26_27,N0_27_27,N3_0_27,N4_10_27,N4_11_28);
-- In matrix 3 adding FA to column 27 
	-- signal N4_12_27 : std_logic;
	-- signal N4_13_28 : std_logic;
	FA899 : full_adder port map (N3_1_27,N3_2_27,N3_3_27,N4_12_27,N4_13_28);
-- In matrix 3 adding FA to column 27 
	-- signal N4_14_27 : std_logic;
	-- signal N4_15_28 : std_logic;
	FA900 : full_adder port map (N3_4_27,N3_5_27,N3_6_27,N4_14_27,N4_15_28);
-- In matrix 3 adding FA to column 28 
	-- signal N4_0_28 : std_logic;
	-- signal N4_1_29 : std_logic;
	FA901 : full_adder port map (N0_14_28,N0_15_28,N0_16_28,N4_0_28,N4_1_29);
-- In matrix 3 adding FA to column 28 
	-- signal N4_2_28 : std_logic;
	-- signal N4_3_29 : std_logic;
	FA902 : full_adder port map (N0_17_28,N0_18_28,N0_19_28,N4_2_28,N4_3_29);
-- In matrix 3 adding FA to column 28 
	-- signal N4_4_28 : std_logic;
	-- signal N4_5_29 : std_logic;
	FA903 : full_adder port map (N0_20_28,N0_21_28,N0_22_28,N4_4_28,N4_5_29);
-- In matrix 3 adding FA to column 28 
	-- signal N4_6_28 : std_logic;
	-- signal N4_7_29 : std_logic;
	FA904 : full_adder port map (N0_23_28,N0_24_28,N0_25_28,N4_6_28,N4_7_29);
-- In matrix 3 adding FA to column 28 
	-- signal N4_8_28 : std_logic;
	-- signal N4_9_29 : std_logic;
	FA905 : full_adder port map (N0_26_28,N0_27_28,N0_28_28,N4_8_28,N4_9_29);
-- In matrix 3 adding FA to column 28 
	-- signal N4_10_28 : std_logic;
	-- signal N4_11_29 : std_logic;
	FA906 : full_adder port map (N3_0_28,N3_1_28,N3_2_28,N4_10_28,N4_11_29);
-- In matrix 3 adding FA to column 28 
	-- signal N4_12_28 : std_logic;
	-- signal N4_13_29 : std_logic;
	FA907 : full_adder port map (N3_3_28,N3_4_28,N3_5_28,N4_12_28,N4_13_29);
-- In matrix 3 adding FA to column 28 
	-- signal N4_14_28 : std_logic;
	-- signal N4_15_29 : std_logic;
	FA908 : full_adder port map (N3_6_28,N3_7_28,N3_8_28,N4_14_28,N4_15_29);
-- In matrix 3 adding FA to column 29 
	-- signal N4_0_29 : std_logic;
	-- signal N4_1_30 : std_logic;
	FA909 : full_adder port map (N0_17_29,N0_18_29,N0_19_29,N4_0_29,N4_1_30);
-- In matrix 3 adding FA to column 29 
	-- signal N4_2_29 : std_logic;
	-- signal N4_3_30 : std_logic;
	FA910 : full_adder port map (N0_20_29,N0_21_29,N0_22_29,N4_2_29,N4_3_30);
-- In matrix 3 adding FA to column 29 
	-- signal N4_4_29 : std_logic;
	-- signal N4_5_30 : std_logic;
	FA911 : full_adder port map (N0_23_29,N0_24_29,N0_25_29,N4_4_29,N4_5_30);
-- In matrix 3 adding FA to column 29 
	-- signal N4_6_29 : std_logic;
	-- signal N4_7_30 : std_logic;
	FA912 : full_adder port map (N0_26_29,N0_27_29,N0_28_29,N4_6_29,N4_7_30);
-- In matrix 3 adding FA to column 29 
	-- signal N4_8_29 : std_logic;
	-- signal N4_9_30 : std_logic;
	FA913 : full_adder port map (N0_29_29,N3_0_29,N3_1_29,N4_8_29,N4_9_30);
-- In matrix 3 adding FA to column 29 
	-- signal N4_10_29 : std_logic;
	-- signal N4_11_30 : std_logic;
	FA914 : full_adder port map (N3_2_29,N3_3_29,N3_4_29,N4_10_29,N4_11_30);
-- In matrix 3 adding FA to column 29 
	-- signal N4_12_29 : std_logic;
	-- signal N4_13_30 : std_logic;
	FA915 : full_adder port map (N3_5_29,N3_6_29,N3_7_29,N4_12_29,N4_13_30);
-- In matrix 3 adding FA to column 29 
	-- signal N4_14_29 : std_logic;
	-- signal N4_15_30 : std_logic;
	FA916 : full_adder port map (N3_8_29,N3_9_29,N3_10_29,N4_14_29,N4_15_30);
-- In matrix 3 adding FA to column 30 
	-- signal N4_0_30 : std_logic;
	-- signal N4_1_31 : std_logic;
	FA917 : full_adder port map (N0_20_30,N0_21_30,N0_22_30,N4_0_30,N4_1_31);
-- In matrix 3 adding FA to column 30 
	-- signal N4_2_30 : std_logic;
	-- signal N4_3_31 : std_logic;
	FA918 : full_adder port map (N0_23_30,N0_24_30,N0_25_30,N4_2_30,N4_3_31);
-- In matrix 3 adding FA to column 30 
	-- signal N4_4_30 : std_logic;
	-- signal N4_5_31 : std_logic;
	FA919 : full_adder port map (N0_26_30,N0_27_30,N0_28_30,N4_4_30,N4_5_31);
-- In matrix 3 adding FA to column 30 
	-- signal N4_6_30 : std_logic;
	-- signal N4_7_31 : std_logic;
	FA920 : full_adder port map (N0_29_30,N0_30_30,N3_0_30,N4_6_30,N4_7_31);
-- In matrix 3 adding FA to column 30 
	-- signal N4_8_30 : std_logic;
	-- signal N4_9_31 : std_logic;
	FA921 : full_adder port map (N3_1_30,N3_2_30,N3_3_30,N4_8_30,N4_9_31);
-- In matrix 3 adding FA to column 30 
	-- signal N4_10_30 : std_logic;
	-- signal N4_11_31 : std_logic;
	FA922 : full_adder port map (N3_4_30,N3_5_30,N3_6_30,N4_10_30,N4_11_31);
-- In matrix 3 adding FA to column 30 
	-- signal N4_12_30 : std_logic;
	-- signal N4_13_31 : std_logic;
	FA923 : full_adder port map (N3_7_30,N3_8_30,N3_9_30,N4_12_30,N4_13_31);
-- In matrix 3 adding FA to column 30 
	-- signal N4_14_30 : std_logic;
	-- signal N4_15_31 : std_logic;
	FA924 : full_adder port map (N3_10_30,N3_11_30,N3_12_30,N4_14_30,N4_15_31);
-- In matrix 3 adding FA to column 31 
	-- signal N4_0_31 : std_logic;
	-- signal N4_1_32 : std_logic;
	FA925 : full_adder port map (N0_23_31,N0_24_31,N0_25_31,N4_0_31,N4_1_32);
-- In matrix 3 adding FA to column 31 
	-- signal N4_2_31 : std_logic;
	-- signal N4_3_32 : std_logic;
	FA926 : full_adder port map (N0_26_31,N0_27_31,N0_28_31,N4_2_31,N4_3_32);
-- In matrix 3 adding FA to column 31 
	-- signal N4_4_31 : std_logic;
	-- signal N4_5_32 : std_logic;
	FA927 : full_adder port map (N0_29_31,N0_30_31,N0_31_31,N4_4_31,N4_5_32);
-- In matrix 3 adding FA to column 31 
	-- signal N4_6_31 : std_logic;
	-- signal N4_7_32 : std_logic;
	FA928 : full_adder port map (N3_0_31,N3_1_31,N3_2_31,N4_6_31,N4_7_32);
-- In matrix 3 adding FA to column 31 
	-- signal N4_8_31 : std_logic;
	-- signal N4_9_32 : std_logic;
	FA929 : full_adder port map (N3_3_31,N3_4_31,N3_5_31,N4_8_31,N4_9_32);
-- In matrix 3 adding FA to column 31 
	-- signal N4_10_31 : std_logic;
	-- signal N4_11_32 : std_logic;
	FA930 : full_adder port map (N3_6_31,N3_7_31,N3_8_31,N4_10_31,N4_11_32);
-- In matrix 3 adding FA to column 31 
	-- signal N4_12_31 : std_logic;
	-- signal N4_13_32 : std_logic;
	FA931 : full_adder port map (N3_9_31,N3_10_31,N3_11_31,N4_12_31,N4_13_32);
-- In matrix 3 adding FA to column 31 
	-- signal N4_14_31 : std_logic;
	-- signal N4_15_32 : std_logic;
	FA932 : full_adder port map (N3_12_31,N3_13_31,N3_14_31,N4_14_31,N4_15_32);
-- In matrix 3 adding FA to column 32 
	-- signal N4_0_32 : std_logic;
	-- signal N4_1_33 : std_logic;
	FA933 : full_adder port map (N0_26_32,N0_27_32,N0_28_32,N4_0_32,N4_1_33);
-- In matrix 3 adding FA to column 32 
	-- signal N4_2_32 : std_logic;
	-- signal N4_3_33 : std_logic;
	FA934 : full_adder port map (N0_29_32,N0_30_32,N0_31_32,N4_2_32,N4_3_33);
-- In matrix 3 adding FA to column 32 
	-- signal N4_4_32 : std_logic;
	-- signal N4_5_33 : std_logic;
	FA935 : full_adder port map (N0_32_32,N3_0_32,N3_1_32,N4_4_32,N4_5_33);
-- In matrix 3 adding FA to column 32 
	-- signal N4_6_32 : std_logic;
	-- signal N4_7_33 : std_logic;
	FA936 : full_adder port map (N3_2_32,N3_3_32,N3_4_32,N4_6_32,N4_7_33);
-- In matrix 3 adding FA to column 32 
	-- signal N4_8_32 : std_logic;
	-- signal N4_9_33 : std_logic;
	FA937 : full_adder port map (N3_5_32,N3_6_32,N3_7_32,N4_8_32,N4_9_33);
-- In matrix 3 adding FA to column 32 
	-- signal N4_10_32 : std_logic;
	-- signal N4_11_33 : std_logic;
	FA938 : full_adder port map (N3_8_32,N3_9_32,N3_10_32,N4_10_32,N4_11_33);
-- In matrix 3 adding FA to column 32 
	-- signal N4_12_32 : std_logic;
	-- signal N4_13_33 : std_logic;
	FA939 : full_adder port map (N3_11_32,N3_12_32,N3_13_32,N4_12_32,N4_13_33);
-- In matrix 3 adding FA to column 32 
	-- signal N4_14_32 : std_logic;
	-- signal N4_15_33 : std_logic;
	FA940 : full_adder port map (N3_14_32,N3_15_32,N3_16_32,N4_14_32,N4_15_33);
-- In matrix 3 adding FA to column 33 
	-- signal N4_0_33 : std_logic;
	-- signal N4_1_34 : std_logic;
	FA941 : full_adder port map (N0_29_33,N0_30_33,N0_31_33,N4_0_33,N4_1_34);
-- In matrix 3 adding FA to column 33 
	-- signal N4_2_33 : std_logic;
	-- signal N4_3_34 : std_logic;
	FA942 : full_adder port map (N0_32_33,N0_33_33,N3_0_33,N4_2_33,N4_3_34);
-- In matrix 3 adding FA to column 33 
	-- signal N4_4_33 : std_logic;
	-- signal N4_5_34 : std_logic;
	FA943 : full_adder port map (N3_1_33,N3_2_33,N3_3_33,N4_4_33,N4_5_34);
-- In matrix 3 adding FA to column 33 
	-- signal N4_6_33 : std_logic;
	-- signal N4_7_34 : std_logic;
	FA944 : full_adder port map (N3_4_33,N3_5_33,N3_6_33,N4_6_33,N4_7_34);
-- In matrix 3 adding FA to column 33 
	-- signal N4_8_33 : std_logic;
	-- signal N4_9_34 : std_logic;
	FA945 : full_adder port map (N3_7_33,N3_8_33,N3_9_33,N4_8_33,N4_9_34);
-- In matrix 3 adding FA to column 33 
	-- signal N4_10_33 : std_logic;
	-- signal N4_11_34 : std_logic;
	FA946 : full_adder port map (N3_10_33,N3_11_33,N3_12_33,N4_10_33,N4_11_34);
-- In matrix 3 adding FA to column 33 
	-- signal N4_12_33 : std_logic;
	-- signal N4_13_34 : std_logic;
	FA947 : full_adder port map (N3_13_33,N3_14_33,N3_15_33,N4_12_33,N4_13_34);
-- In matrix 3 adding FA to column 33 
	-- signal N4_14_33 : std_logic;
	-- signal N4_15_34 : std_logic;
	FA948 : full_adder port map (N3_16_33,N3_17_33,N3_18_33,N4_14_33,N4_15_34);
-- In matrix 3 adding FA to column 34 
	-- signal N4_0_34 : std_logic;
	-- signal N4_1_35 : std_logic;
	FA949 : full_adder port map (N0_32_34,N0_33_34,N0_34_34,N4_0_34,N4_1_35);
-- In matrix 3 adding FA to column 34 
	-- signal N4_2_34 : std_logic;
	-- signal N4_3_35 : std_logic;
	FA950 : full_adder port map (N3_0_34,N3_1_34,N3_2_34,N4_2_34,N4_3_35);
-- In matrix 3 adding FA to column 34 
	-- signal N4_4_34 : std_logic;
	-- signal N4_5_35 : std_logic;
	FA951 : full_adder port map (N3_3_34,N3_4_34,N3_5_34,N4_4_34,N4_5_35);
-- In matrix 3 adding FA to column 34 
	-- signal N4_6_34 : std_logic;
	-- signal N4_7_35 : std_logic;
	FA952 : full_adder port map (N3_6_34,N3_7_34,N3_8_34,N4_6_34,N4_7_35);
-- In matrix 3 adding FA to column 34 
	-- signal N4_8_34 : std_logic;
	-- signal N4_9_35 : std_logic;
	FA953 : full_adder port map (N3_9_34,N3_10_34,N3_11_34,N4_8_34,N4_9_35);
-- In matrix 3 adding FA to column 34 
	-- signal N4_10_34 : std_logic;
	-- signal N4_11_35 : std_logic;
	FA954 : full_adder port map (N3_12_34,N3_13_34,N3_14_34,N4_10_34,N4_11_35);
-- In matrix 3 adding FA to column 34 
	-- signal N4_12_34 : std_logic;
	-- signal N4_13_35 : std_logic;
	FA955 : full_adder port map (N3_15_34,N3_16_34,N3_17_34,N4_12_34,N4_13_35);
-- In matrix 3 adding FA to column 34 
	-- signal N4_14_34 : std_logic;
	-- signal N4_15_35 : std_logic;
	FA956 : full_adder port map (N3_18_34,N3_19_34,N3_20_34,N4_14_34,N4_15_35);
-- In matrix 3 adding FA to column 35 
	-- signal N4_0_35 : std_logic;
	-- signal N4_1_36 : std_logic;
	FA957 : full_adder port map (N0_35_35,N3_0_35,N3_1_35,N4_0_35,N4_1_36);
-- In matrix 3 adding FA to column 35 
	-- signal N4_2_35 : std_logic;
	-- signal N4_3_36 : std_logic;
	FA958 : full_adder port map (N3_2_35,N3_3_35,N3_4_35,N4_2_35,N4_3_36);
-- In matrix 3 adding FA to column 35 
	-- signal N4_4_35 : std_logic;
	-- signal N4_5_36 : std_logic;
	FA959 : full_adder port map (N3_5_35,N3_6_35,N3_7_35,N4_4_35,N4_5_36);
-- In matrix 3 adding FA to column 35 
	-- signal N4_6_35 : std_logic;
	-- signal N4_7_36 : std_logic;
	FA960 : full_adder port map (N3_8_35,N3_9_35,N3_10_35,N4_6_35,N4_7_36);
-- In matrix 3 adding FA to column 35 
	-- signal N4_8_35 : std_logic;
	-- signal N4_9_36 : std_logic;
	FA961 : full_adder port map (N3_11_35,N3_12_35,N3_13_35,N4_8_35,N4_9_36);
-- In matrix 3 adding FA to column 35 
	-- signal N4_10_35 : std_logic;
	-- signal N4_11_36 : std_logic;
	FA962 : full_adder port map (N3_14_35,N3_15_35,N3_16_35,N4_10_35,N4_11_36);
-- In matrix 3 adding FA to column 35 
	-- signal N4_12_35 : std_logic;
	-- signal N4_13_36 : std_logic;
	FA963 : full_adder port map (N3_17_35,N3_18_35,N3_19_35,N4_12_35,N4_13_36);
-- In matrix 3 adding FA to column 35 
	-- signal N4_14_35 : std_logic;
	-- signal N4_15_36 : std_logic;
	FA964 : full_adder port map (N3_20_35,N3_21_35,N3_22_35,N4_14_35,N4_15_36);
-- In matrix 3 adding FA to column 36 
	-- signal N4_0_36 : std_logic;
	-- signal N4_1_37 : std_logic;
	FA965 : full_adder port map (N3_0_36,N3_1_36,N3_2_36,N4_0_36,N4_1_37);
-- In matrix 3 adding FA to column 36 
	-- signal N4_2_36 : std_logic;
	-- signal N4_3_37 : std_logic;
	FA966 : full_adder port map (N3_3_36,N3_4_36,N3_5_36,N4_2_36,N4_3_37);
-- In matrix 3 adding FA to column 36 
	-- signal N4_4_36 : std_logic;
	-- signal N4_5_37 : std_logic;
	FA967 : full_adder port map (N3_6_36,N3_7_36,N3_8_36,N4_4_36,N4_5_37);
-- In matrix 3 adding FA to column 36 
	-- signal N4_6_36 : std_logic;
	-- signal N4_7_37 : std_logic;
	FA968 : full_adder port map (N3_9_36,N3_10_36,N3_11_36,N4_6_36,N4_7_37);
-- In matrix 3 adding FA to column 36 
	-- signal N4_8_36 : std_logic;
	-- signal N4_9_37 : std_logic;
	FA969 : full_adder port map (N3_12_36,N3_13_36,N3_14_36,N4_8_36,N4_9_37);
-- In matrix 3 adding FA to column 36 
	-- signal N4_10_36 : std_logic;
	-- signal N4_11_37 : std_logic;
	FA970 : full_adder port map (N3_15_36,N3_16_36,N3_17_36,N4_10_36,N4_11_37);
-- In matrix 3 adding FA to column 36 
	-- signal N4_12_36 : std_logic;
	-- signal N4_13_37 : std_logic;
	FA971 : full_adder port map (N3_18_36,N3_19_36,N3_20_36,N4_12_36,N4_13_37);
-- In matrix 3 adding FA to column 36 
	-- signal N4_14_36 : std_logic;
	-- signal N4_15_37 : std_logic;
	FA972 : full_adder port map (N3_21_36,N3_22_36,N3_23_36,N4_14_36,N4_15_37);
-- In matrix 3 adding FA to column 37 
	-- signal N4_0_37 : std_logic;
	-- signal N4_1_38 : std_logic;
	FA973 : full_adder port map (N3_0_37,N3_1_37,N3_2_37,N4_0_37,N4_1_38);
-- In matrix 3 adding FA to column 37 
	-- signal N4_2_37 : std_logic;
	-- signal N4_3_38 : std_logic;
	FA974 : full_adder port map (N3_3_37,N3_4_37,N3_5_37,N4_2_37,N4_3_38);
-- In matrix 3 adding FA to column 37 
	-- signal N4_4_37 : std_logic;
	-- signal N4_5_38 : std_logic;
	FA975 : full_adder port map (N3_6_37,N3_7_37,N3_8_37,N4_4_37,N4_5_38);
-- In matrix 3 adding FA to column 37 
	-- signal N4_6_37 : std_logic;
	-- signal N4_7_38 : std_logic;
	FA976 : full_adder port map (N3_9_37,N3_10_37,N3_11_37,N4_6_37,N4_7_38);
-- In matrix 3 adding FA to column 37 
	-- signal N4_8_37 : std_logic;
	-- signal N4_9_38 : std_logic;
	FA977 : full_adder port map (N3_12_37,N3_13_37,N3_14_37,N4_8_37,N4_9_38);
-- In matrix 3 adding FA to column 37 
	-- signal N4_10_37 : std_logic;
	-- signal N4_11_38 : std_logic;
	FA978 : full_adder port map (N3_15_37,N3_16_37,N3_17_37,N4_10_37,N4_11_38);
-- In matrix 3 adding FA to column 37 
	-- signal N4_12_37 : std_logic;
	-- signal N4_13_38 : std_logic;
	FA979 : full_adder port map (N3_18_37,N3_19_37,N3_20_37,N4_12_37,N4_13_38);
-- In matrix 3 adding FA to column 37 
	-- signal N4_14_37 : std_logic;
	-- signal N4_15_38 : std_logic;
	FA980 : full_adder port map (N3_21_37,N3_22_37,N3_23_37,N4_14_37,N4_15_38);
-- In matrix 3 adding FA to column 38 
	-- signal N4_0_38 : std_logic;
	-- signal N4_1_39 : std_logic;
	FA981 : full_adder port map (N3_0_38,N3_1_38,N3_2_38,N4_0_38,N4_1_39);
-- In matrix 3 adding FA to column 38 
	-- signal N4_2_38 : std_logic;
	-- signal N4_3_39 : std_logic;
	FA982 : full_adder port map (N3_3_38,N3_4_38,N3_5_38,N4_2_38,N4_3_39);
-- In matrix 3 adding FA to column 38 
	-- signal N4_4_38 : std_logic;
	-- signal N4_5_39 : std_logic;
	FA983 : full_adder port map (N3_6_38,N3_7_38,N3_8_38,N4_4_38,N4_5_39);
-- In matrix 3 adding FA to column 38 
	-- signal N4_6_38 : std_logic;
	-- signal N4_7_39 : std_logic;
	FA984 : full_adder port map (N3_9_38,N3_10_38,N3_11_38,N4_6_38,N4_7_39);
-- In matrix 3 adding FA to column 38 
	-- signal N4_8_38 : std_logic;
	-- signal N4_9_39 : std_logic;
	FA985 : full_adder port map (N3_12_38,N3_13_38,N3_14_38,N4_8_38,N4_9_39);
-- In matrix 3 adding FA to column 38 
	-- signal N4_10_38 : std_logic;
	-- signal N4_11_39 : std_logic;
	FA986 : full_adder port map (N3_15_38,N3_16_38,N3_17_38,N4_10_38,N4_11_39);
-- In matrix 3 adding FA to column 38 
	-- signal N4_12_38 : std_logic;
	-- signal N4_13_39 : std_logic;
	FA987 : full_adder port map (N3_18_38,N3_19_38,N3_20_38,N4_12_38,N4_13_39);
-- In matrix 3 adding FA to column 38 
	-- signal N4_14_38 : std_logic;
	-- signal N4_15_39 : std_logic;
	FA988 : full_adder port map (N3_21_38,N3_22_38,N3_23_38,N4_14_38,N4_15_39);
-- In matrix 3 adding FA to column 39 
	-- signal N4_0_39 : std_logic;
	-- signal N4_1_40 : std_logic;
	FA989 : full_adder port map (N3_0_39,N3_1_39,N3_2_39,N4_0_39,N4_1_40);
-- In matrix 3 adding FA to column 39 
	-- signal N4_2_39 : std_logic;
	-- signal N4_3_40 : std_logic;
	FA990 : full_adder port map (N3_3_39,N3_4_39,N3_5_39,N4_2_39,N4_3_40);
-- In matrix 3 adding FA to column 39 
	-- signal N4_4_39 : std_logic;
	-- signal N4_5_40 : std_logic;
	FA991 : full_adder port map (N3_6_39,N3_7_39,N3_8_39,N4_4_39,N4_5_40);
-- In matrix 3 adding FA to column 39 
	-- signal N4_6_39 : std_logic;
	-- signal N4_7_40 : std_logic;
	FA992 : full_adder port map (N3_9_39,N3_10_39,N3_11_39,N4_6_39,N4_7_40);
-- In matrix 3 adding FA to column 39 
	-- signal N4_8_39 : std_logic;
	-- signal N4_9_40 : std_logic;
	FA993 : full_adder port map (N3_12_39,N3_13_39,N3_14_39,N4_8_39,N4_9_40);
-- In matrix 3 adding FA to column 39 
	-- signal N4_10_39 : std_logic;
	-- signal N4_11_40 : std_logic;
	FA994 : full_adder port map (N3_15_39,N3_16_39,N3_17_39,N4_10_39,N4_11_40);
-- In matrix 3 adding FA to column 39 
	-- signal N4_12_39 : std_logic;
	-- signal N4_13_40 : std_logic;
	FA995 : full_adder port map (N3_18_39,N3_19_39,N3_20_39,N4_12_39,N4_13_40);
-- In matrix 3 adding FA to column 39 
	-- signal N4_14_39 : std_logic;
	-- signal N4_15_40 : std_logic;
	FA996 : full_adder port map (N3_21_39,N3_22_39,N3_23_39,N4_14_39,N4_15_40);
-- In matrix 3 adding FA to column 40 
	-- signal N4_0_40 : std_logic;
	-- signal N4_1_41 : std_logic;
	FA997 : full_adder port map (N3_0_40,N3_1_40,N3_2_40,N4_0_40,N4_1_41);
-- In matrix 3 adding FA to column 40 
	-- signal N4_2_40 : std_logic;
	-- signal N4_3_41 : std_logic;
	FA998 : full_adder port map (N3_3_40,N3_4_40,N3_5_40,N4_2_40,N4_3_41);
-- In matrix 3 adding FA to column 40 
	-- signal N4_4_40 : std_logic;
	-- signal N4_5_41 : std_logic;
	FA999 : full_adder port map (N3_6_40,N3_7_40,N3_8_40,N4_4_40,N4_5_41);
-- In matrix 3 adding FA to column 40 
	-- signal N4_6_40 : std_logic;
	-- signal N4_7_41 : std_logic;
	FA1000 : full_adder port map (N3_9_40,N3_10_40,N3_11_40,N4_6_40,N4_7_41);
-- In matrix 3 adding FA to column 40 
	-- signal N4_8_40 : std_logic;
	-- signal N4_9_41 : std_logic;
	FA1001 : full_adder port map (N3_12_40,N3_13_40,N3_14_40,N4_8_40,N4_9_41);
-- In matrix 3 adding FA to column 40 
	-- signal N4_10_40 : std_logic;
	-- signal N4_11_41 : std_logic;
	FA1002 : full_adder port map (N3_15_40,N3_16_40,N3_17_40,N4_10_40,N4_11_41);
-- In matrix 3 adding FA to column 40 
	-- signal N4_12_40 : std_logic;
	-- signal N4_13_41 : std_logic;
	FA1003 : full_adder port map (N3_18_40,N3_19_40,N3_20_40,N4_12_40,N4_13_41);
-- In matrix 3 adding FA to column 40 
	-- signal N4_14_40 : std_logic;
	-- signal N4_15_41 : std_logic;
	FA1004 : full_adder port map (N3_21_40,N3_22_40,N3_23_40,N4_14_40,N4_15_41);
-- In matrix 3 adding FA to column 41 
	-- signal N4_0_41 : std_logic;
	-- signal N4_1_42 : std_logic;
	FA1005 : full_adder port map (N3_0_41,N3_1_41,N3_2_41,N4_0_41,N4_1_42);
-- In matrix 3 adding FA to column 41 
	-- signal N4_2_41 : std_logic;
	-- signal N4_3_42 : std_logic;
	FA1006 : full_adder port map (N3_3_41,N3_4_41,N3_5_41,N4_2_41,N4_3_42);
-- In matrix 3 adding FA to column 41 
	-- signal N4_4_41 : std_logic;
	-- signal N4_5_42 : std_logic;
	FA1007 : full_adder port map (N3_6_41,N3_7_41,N3_8_41,N4_4_41,N4_5_42);
-- In matrix 3 adding FA to column 41 
	-- signal N4_6_41 : std_logic;
	-- signal N4_7_42 : std_logic;
	FA1008 : full_adder port map (N3_9_41,N3_10_41,N3_11_41,N4_6_41,N4_7_42);
-- In matrix 3 adding FA to column 41 
	-- signal N4_8_41 : std_logic;
	-- signal N4_9_42 : std_logic;
	FA1009 : full_adder port map (N3_12_41,N3_13_41,N3_14_41,N4_8_41,N4_9_42);
-- In matrix 3 adding FA to column 41 
	-- signal N4_10_41 : std_logic;
	-- signal N4_11_42 : std_logic;
	FA1010 : full_adder port map (N3_15_41,N3_16_41,N3_17_41,N4_10_41,N4_11_42);
-- In matrix 3 adding FA to column 41 
	-- signal N4_12_41 : std_logic;
	-- signal N4_13_42 : std_logic;
	FA1011 : full_adder port map (N3_18_41,N3_19_41,N3_20_41,N4_12_41,N4_13_42);
-- In matrix 3 adding FA to column 41 
	-- signal N4_14_41 : std_logic;
	-- signal N4_15_42 : std_logic;
	FA1012 : full_adder port map (N3_21_41,N3_22_41,N3_23_41,N4_14_41,N4_15_42);
-- In matrix 3 adding FA to column 42 
	-- signal N4_0_42 : std_logic;
	-- signal N4_1_43 : std_logic;
	FA1013 : full_adder port map (N3_0_42,N3_1_42,N3_2_42,N4_0_42,N4_1_43);
-- In matrix 3 adding FA to column 42 
	-- signal N4_2_42 : std_logic;
	-- signal N4_3_43 : std_logic;
	FA1014 : full_adder port map (N3_3_42,N3_4_42,N3_5_42,N4_2_42,N4_3_43);
-- In matrix 3 adding FA to column 42 
	-- signal N4_4_42 : std_logic;
	-- signal N4_5_43 : std_logic;
	FA1015 : full_adder port map (N3_6_42,N3_7_42,N3_8_42,N4_4_42,N4_5_43);
-- In matrix 3 adding FA to column 42 
	-- signal N4_6_42 : std_logic;
	-- signal N4_7_43 : std_logic;
	FA1016 : full_adder port map (N3_9_42,N3_10_42,N3_11_42,N4_6_42,N4_7_43);
-- In matrix 3 adding FA to column 42 
	-- signal N4_8_42 : std_logic;
	-- signal N4_9_43 : std_logic;
	FA1017 : full_adder port map (N3_12_42,N3_13_42,N3_14_42,N4_8_42,N4_9_43);
-- In matrix 3 adding FA to column 42 
	-- signal N4_10_42 : std_logic;
	-- signal N4_11_43 : std_logic;
	FA1018 : full_adder port map (N3_15_42,N3_16_42,N3_17_42,N4_10_42,N4_11_43);
-- In matrix 3 adding FA to column 42 
	-- signal N4_12_42 : std_logic;
	-- signal N4_13_43 : std_logic;
	FA1019 : full_adder port map (N3_18_42,N3_19_42,N3_20_42,N4_12_42,N4_13_43);
-- In matrix 3 adding FA to column 42 
	-- signal N4_14_42 : std_logic;
	-- signal N4_15_43 : std_logic;
	FA1020 : full_adder port map (N3_21_42,N3_22_42,N3_23_42,N4_14_42,N4_15_43);
-- In matrix 3 adding FA to column 43 
	-- signal N4_0_43 : std_logic;
	-- signal N4_1_44 : std_logic;
	FA1021 : full_adder port map (N3_0_43,N3_1_43,N3_2_43,N4_0_43,N4_1_44);
-- In matrix 3 adding FA to column 43 
	-- signal N4_2_43 : std_logic;
	-- signal N4_3_44 : std_logic;
	FA1022 : full_adder port map (N3_3_43,N3_4_43,N3_5_43,N4_2_43,N4_3_44);
-- In matrix 3 adding FA to column 43 
	-- signal N4_4_43 : std_logic;
	-- signal N4_5_44 : std_logic;
	FA1023 : full_adder port map (N3_6_43,N3_7_43,N3_8_43,N4_4_43,N4_5_44);
-- In matrix 3 adding FA to column 43 
	-- signal N4_6_43 : std_logic;
	-- signal N4_7_44 : std_logic;
	FA1024 : full_adder port map (N3_9_43,N3_10_43,N3_11_43,N4_6_43,N4_7_44);
-- In matrix 3 adding FA to column 43 
	-- signal N4_8_43 : std_logic;
	-- signal N4_9_44 : std_logic;
	FA1025 : full_adder port map (N3_12_43,N3_13_43,N3_14_43,N4_8_43,N4_9_44);
-- In matrix 3 adding FA to column 43 
	-- signal N4_10_43 : std_logic;
	-- signal N4_11_44 : std_logic;
	FA1026 : full_adder port map (N3_15_43,N3_16_43,N3_17_43,N4_10_43,N4_11_44);
-- In matrix 3 adding FA to column 43 
	-- signal N4_12_43 : std_logic;
	-- signal N4_13_44 : std_logic;
	FA1027 : full_adder port map (N3_18_43,N3_19_43,N3_20_43,N4_12_43,N4_13_44);
-- In matrix 3 adding FA to column 43 
	-- signal N4_14_43 : std_logic;
	-- signal N4_15_44 : std_logic;
	FA1028 : full_adder port map (N3_21_43,N3_22_43,N3_23_43,N4_14_43,N4_15_44);
-- In matrix 3 adding FA to column 44 
	-- signal N4_0_44 : std_logic;
	-- signal N4_1_45 : std_logic;
	FA1029 : full_adder port map (N3_0_44,N3_1_44,N3_2_44,N4_0_44,N4_1_45);
-- In matrix 3 adding FA to column 44 
	-- signal N4_2_44 : std_logic;
	-- signal N4_3_45 : std_logic;
	FA1030 : full_adder port map (N3_3_44,N3_4_44,N3_5_44,N4_2_44,N4_3_45);
-- In matrix 3 adding FA to column 44 
	-- signal N4_4_44 : std_logic;
	-- signal N4_5_45 : std_logic;
	FA1031 : full_adder port map (N3_6_44,N3_7_44,N3_8_44,N4_4_44,N4_5_45);
-- In matrix 3 adding FA to column 44 
	-- signal N4_6_44 : std_logic;
	-- signal N4_7_45 : std_logic;
	FA1032 : full_adder port map (N3_9_44,N3_10_44,N3_11_44,N4_6_44,N4_7_45);
-- In matrix 3 adding FA to column 44 
	-- signal N4_8_44 : std_logic;
	-- signal N4_9_45 : std_logic;
	FA1033 : full_adder port map (N3_12_44,N3_13_44,N3_14_44,N4_8_44,N4_9_45);
-- In matrix 3 adding FA to column 44 
	-- signal N4_10_44 : std_logic;
	-- signal N4_11_45 : std_logic;
	FA1034 : full_adder port map (N3_15_44,N3_16_44,N3_17_44,N4_10_44,N4_11_45);
-- In matrix 3 adding FA to column 44 
	-- signal N4_12_44 : std_logic;
	-- signal N4_13_45 : std_logic;
	FA1035 : full_adder port map (N3_18_44,N3_19_44,N3_20_44,N4_12_44,N4_13_45);
-- In matrix 3 adding FA to column 44 
	-- signal N4_14_44 : std_logic;
	-- signal N4_15_45 : std_logic;
	FA1036 : full_adder port map (N3_21_44,N3_22_44,N3_23_44,N4_14_44,N4_15_45);
-- In matrix 3 adding FA to column 45 
	-- signal N4_0_45 : std_logic;
	-- signal N4_1_46 : std_logic;
	FA1037 : full_adder port map (N3_0_45,N3_1_45,N3_2_45,N4_0_45,N4_1_46);
-- In matrix 3 adding FA to column 45 
	-- signal N4_2_45 : std_logic;
	-- signal N4_3_46 : std_logic;
	FA1038 : full_adder port map (N3_3_45,N3_4_45,N3_5_45,N4_2_45,N4_3_46);
-- In matrix 3 adding FA to column 45 
	-- signal N4_4_45 : std_logic;
	-- signal N4_5_46 : std_logic;
	FA1039 : full_adder port map (N3_6_45,N3_7_45,N3_8_45,N4_4_45,N4_5_46);
-- In matrix 3 adding FA to column 45 
	-- signal N4_6_45 : std_logic;
	-- signal N4_7_46 : std_logic;
	FA1040 : full_adder port map (N3_9_45,N3_10_45,N3_11_45,N4_6_45,N4_7_46);
-- In matrix 3 adding FA to column 45 
	-- signal N4_8_45 : std_logic;
	-- signal N4_9_46 : std_logic;
	FA1041 : full_adder port map (N3_12_45,N3_13_45,N3_14_45,N4_8_45,N4_9_46);
-- In matrix 3 adding FA to column 45 
	-- signal N4_10_45 : std_logic;
	-- signal N4_11_46 : std_logic;
	FA1042 : full_adder port map (N3_15_45,N3_16_45,N3_17_45,N4_10_45,N4_11_46);
-- In matrix 3 adding FA to column 45 
	-- signal N4_12_45 : std_logic;
	-- signal N4_13_46 : std_logic;
	FA1043 : full_adder port map (N3_18_45,N3_19_45,N3_20_45,N4_12_45,N4_13_46);
-- In matrix 3 adding FA to column 45 
	-- signal N4_14_45 : std_logic;
	-- signal N4_15_46 : std_logic;
	FA1044 : full_adder port map (N3_21_45,N3_22_45,N3_23_45,N4_14_45,N4_15_46);
-- In matrix 3 adding FA to column 46 
	-- signal N4_0_46 : std_logic;
	-- signal N4_1_47 : std_logic;
	FA1045 : full_adder port map (N3_0_46,N3_1_46,N3_2_46,N4_0_46,N4_1_47);
-- In matrix 3 adding FA to column 46 
	-- signal N4_2_46 : std_logic;
	-- signal N4_3_47 : std_logic;
	FA1046 : full_adder port map (N3_3_46,N3_4_46,N3_5_46,N4_2_46,N4_3_47);
-- In matrix 3 adding FA to column 46 
	-- signal N4_4_46 : std_logic;
	-- signal N4_5_47 : std_logic;
	FA1047 : full_adder port map (N3_6_46,N3_7_46,N3_8_46,N4_4_46,N4_5_47);
-- In matrix 3 adding FA to column 46 
	-- signal N4_6_46 : std_logic;
	-- signal N4_7_47 : std_logic;
	FA1048 : full_adder port map (N3_9_46,N3_10_46,N3_11_46,N4_6_46,N4_7_47);
-- In matrix 3 adding FA to column 46 
	-- signal N4_8_46 : std_logic;
	-- signal N4_9_47 : std_logic;
	FA1049 : full_adder port map (N3_12_46,N3_13_46,N3_14_46,N4_8_46,N4_9_47);
-- In matrix 3 adding FA to column 46 
	-- signal N4_10_46 : std_logic;
	-- signal N4_11_47 : std_logic;
	FA1050 : full_adder port map (N3_15_46,N3_16_46,N3_17_46,N4_10_46,N4_11_47);
-- In matrix 3 adding FA to column 46 
	-- signal N4_12_46 : std_logic;
	-- signal N4_13_47 : std_logic;
	FA1051 : full_adder port map (N3_18_46,N3_19_46,N3_20_46,N4_12_46,N4_13_47);
-- In matrix 3 adding FA to column 46 
	-- signal N4_14_46 : std_logic;
	-- signal N4_15_47 : std_logic;
	FA1052 : full_adder port map (N3_21_46,N3_22_46,N3_23_46,N4_14_46,N4_15_47);
-- In matrix 3 adding FA to column 47 
	-- signal N4_0_47 : std_logic;
	-- signal N4_1_48 : std_logic;
	FA1053 : full_adder port map (N3_0_47,N3_1_47,N3_2_47,N4_0_47,N4_1_48);
-- In matrix 3 adding FA to column 47 
	-- signal N4_2_47 : std_logic;
	-- signal N4_3_48 : std_logic;
	FA1054 : full_adder port map (N3_3_47,N3_4_47,N3_5_47,N4_2_47,N4_3_48);
-- In matrix 3 adding FA to column 47 
	-- signal N4_4_47 : std_logic;
	-- signal N4_5_48 : std_logic;
	FA1055 : full_adder port map (N3_6_47,N3_7_47,N3_8_47,N4_4_47,N4_5_48);
-- In matrix 3 adding FA to column 47 
	-- signal N4_6_47 : std_logic;
	-- signal N4_7_48 : std_logic;
	FA1056 : full_adder port map (N3_9_47,N3_10_47,N3_11_47,N4_6_47,N4_7_48);
-- In matrix 3 adding FA to column 47 
	-- signal N4_8_47 : std_logic;
	-- signal N4_9_48 : std_logic;
	FA1057 : full_adder port map (N3_12_47,N3_13_47,N3_14_47,N4_8_47,N4_9_48);
-- In matrix 3 adding FA to column 47 
	-- signal N4_10_47 : std_logic;
	-- signal N4_11_48 : std_logic;
	FA1058 : full_adder port map (N3_15_47,N3_16_47,N3_17_47,N4_10_47,N4_11_48);
-- In matrix 3 adding FA to column 47 
	-- signal N4_12_47 : std_logic;
	-- signal N4_13_48 : std_logic;
	FA1059 : full_adder port map (N3_18_47,N3_19_47,N3_20_47,N4_12_47,N4_13_48);
-- In matrix 3 adding FA to column 47 
	-- signal N4_14_47 : std_logic;
	-- signal N4_15_48 : std_logic;
	FA1060 : full_adder port map (N3_21_47,N3_22_47,N3_23_47,N4_14_47,N4_15_48);
-- In matrix 3 adding FA to column 48 
	-- signal N4_0_48 : std_logic;
	-- signal N4_1_49 : std_logic;
	FA1061 : full_adder port map (N3_0_48,N3_1_48,N3_2_48,N4_0_48,N4_1_49);
-- In matrix 3 adding FA to column 48 
	-- signal N4_2_48 : std_logic;
	-- signal N4_3_49 : std_logic;
	FA1062 : full_adder port map (N3_3_48,N3_4_48,N3_5_48,N4_2_48,N4_3_49);
-- In matrix 3 adding FA to column 48 
	-- signal N4_4_48 : std_logic;
	-- signal N4_5_49 : std_logic;
	FA1063 : full_adder port map (N3_6_48,N3_7_48,N3_8_48,N4_4_48,N4_5_49);
-- In matrix 3 adding FA to column 48 
	-- signal N4_6_48 : std_logic;
	-- signal N4_7_49 : std_logic;
	FA1064 : full_adder port map (N3_9_48,N3_10_48,N3_11_48,N4_6_48,N4_7_49);
-- In matrix 3 adding FA to column 48 
	-- signal N4_8_48 : std_logic;
	-- signal N4_9_49 : std_logic;
	FA1065 : full_adder port map (N3_12_48,N3_13_48,N3_14_48,N4_8_48,N4_9_49);
-- In matrix 3 adding FA to column 48 
	-- signal N4_10_48 : std_logic;
	-- signal N4_11_49 : std_logic;
	FA1066 : full_adder port map (N3_15_48,N3_16_48,N3_17_48,N4_10_48,N4_11_49);
-- In matrix 3 adding FA to column 48 
	-- signal N4_12_48 : std_logic;
	-- signal N4_13_49 : std_logic;
	FA1067 : full_adder port map (N3_18_48,N3_19_48,N3_20_48,N4_12_48,N4_13_49);
-- In matrix 3 adding FA to column 48 
	-- signal N4_14_48 : std_logic;
	-- signal N4_15_49 : std_logic;
	FA1068 : full_adder port map (N3_21_48,N3_22_48,N3_23_48,N4_14_48,N4_15_49);
-- In matrix 3 adding FA to column 49 
	-- signal N4_0_49 : std_logic;
	-- signal N4_1_50 : std_logic;
	FA1069 : full_adder port map (N3_0_49,N3_1_49,N3_2_49,N4_0_49,N4_1_50);
-- In matrix 3 adding FA to column 49 
	-- signal N4_2_49 : std_logic;
	-- signal N4_3_50 : std_logic;
	FA1070 : full_adder port map (N3_3_49,N3_4_49,N3_5_49,N4_2_49,N4_3_50);
-- In matrix 3 adding FA to column 49 
	-- signal N4_4_49 : std_logic;
	-- signal N4_5_50 : std_logic;
	FA1071 : full_adder port map (N3_6_49,N3_7_49,N3_8_49,N4_4_49,N4_5_50);
-- In matrix 3 adding FA to column 49 
	-- signal N4_6_49 : std_logic;
	-- signal N4_7_50 : std_logic;
	FA1072 : full_adder port map (N3_9_49,N3_10_49,N3_11_49,N4_6_49,N4_7_50);
-- In matrix 3 adding FA to column 49 
	-- signal N4_8_49 : std_logic;
	-- signal N4_9_50 : std_logic;
	FA1073 : full_adder port map (N3_12_49,N3_13_49,N3_14_49,N4_8_49,N4_9_50);
-- In matrix 3 adding FA to column 49 
	-- signal N4_10_49 : std_logic;
	-- signal N4_11_50 : std_logic;
	FA1074 : full_adder port map (N3_15_49,N3_16_49,N3_17_49,N4_10_49,N4_11_50);
-- In matrix 3 adding FA to column 49 
	-- signal N4_12_49 : std_logic;
	-- signal N4_13_50 : std_logic;
	FA1075 : full_adder port map (N3_18_49,N3_19_49,N3_20_49,N4_12_49,N4_13_50);
-- In matrix 3 adding FA to column 49 
	-- signal N4_14_49 : std_logic;
	-- signal N4_15_50 : std_logic;
	FA1076 : full_adder port map (N3_21_49,N3_22_49,N3_23_49,N4_14_49,N4_15_50);
-- In matrix 3 adding FA to column 50 
	-- signal N4_0_50 : std_logic;
	-- signal N4_1_51 : std_logic;
	FA1077 : full_adder port map (N3_0_50,N3_1_50,N3_2_50,N4_0_50,N4_1_51);
-- In matrix 3 adding FA to column 50 
	-- signal N4_2_50 : std_logic;
	-- signal N4_3_51 : std_logic;
	FA1078 : full_adder port map (N3_3_50,N3_4_50,N3_5_50,N4_2_50,N4_3_51);
-- In matrix 3 adding FA to column 50 
	-- signal N4_4_50 : std_logic;
	-- signal N4_5_51 : std_logic;
	FA1079 : full_adder port map (N3_6_50,N3_7_50,N3_8_50,N4_4_50,N4_5_51);
-- In matrix 3 adding FA to column 50 
	-- signal N4_6_50 : std_logic;
	-- signal N4_7_51 : std_logic;
	FA1080 : full_adder port map (N3_9_50,N3_10_50,N3_11_50,N4_6_50,N4_7_51);
-- In matrix 3 adding FA to column 50 
	-- signal N4_8_50 : std_logic;
	-- signal N4_9_51 : std_logic;
	FA1081 : full_adder port map (N3_12_50,N3_13_50,N3_14_50,N4_8_50,N4_9_51);
-- In matrix 3 adding FA to column 50 
	-- signal N4_10_50 : std_logic;
	-- signal N4_11_51 : std_logic;
	FA1082 : full_adder port map (N3_15_50,N3_16_50,N3_17_50,N4_10_50,N4_11_51);
-- In matrix 3 adding FA to column 50 
	-- signal N4_12_50 : std_logic;
	-- signal N4_13_51 : std_logic;
	FA1083 : full_adder port map (N3_18_50,N3_19_50,N3_20_50,N4_12_50,N4_13_51);
-- In matrix 3 adding FA to column 50 
	-- signal N4_14_50 : std_logic;
	-- signal N4_15_51 : std_logic;
	FA1084 : full_adder port map (N3_21_50,N3_22_50,N3_23_50,N4_14_50,N4_15_51);
-- In matrix 3 adding FA to column 51 
	-- signal N4_0_51 : std_logic;
	-- signal N4_1_52 : std_logic;
	FA1085 : full_adder port map (N3_0_51,N3_1_51,N3_2_51,N4_0_51,N4_1_52);
-- In matrix 3 adding FA to column 51 
	-- signal N4_2_51 : std_logic;
	-- signal N4_3_52 : std_logic;
	FA1086 : full_adder port map (N3_3_51,N3_4_51,N3_5_51,N4_2_51,N4_3_52);
-- In matrix 3 adding FA to column 51 
	-- signal N4_4_51 : std_logic;
	-- signal N4_5_52 : std_logic;
	FA1087 : full_adder port map (N3_6_51,N3_7_51,N3_8_51,N4_4_51,N4_5_52);
-- In matrix 3 adding FA to column 51 
	-- signal N4_6_51 : std_logic;
	-- signal N4_7_52 : std_logic;
	FA1088 : full_adder port map (N3_9_51,N3_10_51,N3_11_51,N4_6_51,N4_7_52);
-- In matrix 3 adding FA to column 51 
	-- signal N4_8_51 : std_logic;
	-- signal N4_9_52 : std_logic;
	FA1089 : full_adder port map (N3_12_51,N3_13_51,N3_14_51,N4_8_51,N4_9_52);
-- In matrix 3 adding FA to column 51 
	-- signal N4_10_51 : std_logic;
	-- signal N4_11_52 : std_logic;
	FA1090 : full_adder port map (N3_15_51,N3_16_51,N3_17_51,N4_10_51,N4_11_52);
-- In matrix 3 adding FA to column 51 
	-- signal N4_12_51 : std_logic;
	-- signal N4_13_52 : std_logic;
	FA1091 : full_adder port map (N3_18_51,N3_19_51,N3_20_51,N4_12_51,N4_13_52);
-- In matrix 3 adding FA to column 51 
	-- signal N4_14_51 : std_logic;
	-- signal N4_15_52 : std_logic;
	FA1092 : full_adder port map (N3_21_51,N3_22_51,N3_23_51,N4_14_51,N4_15_52);
-- In matrix 3 adding FA to column 52 
	-- signal N4_0_52 : std_logic;
	-- signal N4_1_53 : std_logic;
	FA1093 : full_adder port map (N3_0_52,N3_1_52,N3_2_52,N4_0_52,N4_1_53);
-- In matrix 3 adding FA to column 52 
	-- signal N4_2_52 : std_logic;
	-- signal N4_3_53 : std_logic;
	FA1094 : full_adder port map (N3_3_52,N3_4_52,N3_5_52,N4_2_52,N4_3_53);
-- In matrix 3 adding FA to column 52 
	-- signal N4_4_52 : std_logic;
	-- signal N4_5_53 : std_logic;
	FA1095 : full_adder port map (N3_6_52,N3_7_52,N3_8_52,N4_4_52,N4_5_53);
-- In matrix 3 adding FA to column 52 
	-- signal N4_6_52 : std_logic;
	-- signal N4_7_53 : std_logic;
	FA1096 : full_adder port map (N3_9_52,N3_10_52,N3_11_52,N4_6_52,N4_7_53);
-- In matrix 3 adding FA to column 52 
	-- signal N4_8_52 : std_logic;
	-- signal N4_9_53 : std_logic;
	FA1097 : full_adder port map (N3_12_52,N3_13_52,N3_14_52,N4_8_52,N4_9_53);
-- In matrix 3 adding FA to column 52 
	-- signal N4_10_52 : std_logic;
	-- signal N4_11_53 : std_logic;
	FA1098 : full_adder port map (N3_15_52,N3_16_52,N3_17_52,N4_10_52,N4_11_53);
-- In matrix 3 adding FA to column 52 
	-- signal N4_12_52 : std_logic;
	-- signal N4_13_53 : std_logic;
	FA1099 : full_adder port map (N3_18_52,N3_19_52,N3_20_52,N4_12_52,N4_13_53);
-- In matrix 3 adding FA to column 52 
	-- signal N4_14_52 : std_logic;
	-- signal N4_15_53 : std_logic;
	FA1100 : full_adder port map (N3_21_52,N3_22_52,N3_23_52,N4_14_52,N4_15_53);
-- In matrix 3 adding FA to column 53 
	-- signal N4_0_53 : std_logic;
	-- signal N4_1_54 : std_logic;
	FA1101 : full_adder port map (N3_0_53,N3_1_53,N3_2_53,N4_0_53,N4_1_54);
-- In matrix 3 adding FA to column 53 
	-- signal N4_2_53 : std_logic;
	-- signal N4_3_54 : std_logic;
	FA1102 : full_adder port map (N3_3_53,N3_4_53,N3_5_53,N4_2_53,N4_3_54);
-- In matrix 3 adding FA to column 53 
	-- signal N4_4_53 : std_logic;
	-- signal N4_5_54 : std_logic;
	FA1103 : full_adder port map (N3_6_53,N3_7_53,N3_8_53,N4_4_53,N4_5_54);
-- In matrix 3 adding FA to column 53 
	-- signal N4_6_53 : std_logic;
	-- signal N4_7_54 : std_logic;
	FA1104 : full_adder port map (N3_9_53,N3_10_53,N3_11_53,N4_6_53,N4_7_54);
-- In matrix 3 adding FA to column 53 
	-- signal N4_8_53 : std_logic;
	-- signal N4_9_54 : std_logic;
	FA1105 : full_adder port map (N3_12_53,N3_13_53,N3_14_53,N4_8_53,N4_9_54);
-- In matrix 3 adding FA to column 53 
	-- signal N4_10_53 : std_logic;
	-- signal N4_11_54 : std_logic;
	FA1106 : full_adder port map (N3_15_53,N3_16_53,N3_17_53,N4_10_53,N4_11_54);
-- In matrix 3 adding FA to column 53 
	-- signal N4_12_53 : std_logic;
	-- signal N4_13_54 : std_logic;
	FA1107 : full_adder port map (N3_18_53,N3_19_53,N3_20_53,N4_12_53,N4_13_54);
-- In matrix 3 adding FA to column 53 
	-- signal N4_14_53 : std_logic;
	-- signal N4_15_54 : std_logic;
	FA1108 : full_adder port map (N3_21_53,N3_22_53,N3_23_53,N4_14_53,N4_15_54);
-- In matrix 3 adding FA to column 54 
	-- signal N4_0_54 : std_logic;
	-- signal N4_1_55 : std_logic;
	FA1109 : full_adder port map (N3_0_54,N3_1_54,N3_2_54,N4_0_54,N4_1_55);
-- In matrix 3 adding FA to column 54 
	-- signal N4_2_54 : std_logic;
	-- signal N4_3_55 : std_logic;
	FA1110 : full_adder port map (N3_3_54,N3_4_54,N3_5_54,N4_2_54,N4_3_55);
-- In matrix 3 adding FA to column 54 
	-- signal N4_4_54 : std_logic;
	-- signal N4_5_55 : std_logic;
	FA1111 : full_adder port map (N3_6_54,N3_7_54,N3_8_54,N4_4_54,N4_5_55);
-- In matrix 3 adding FA to column 54 
	-- signal N4_6_54 : std_logic;
	-- signal N4_7_55 : std_logic;
	FA1112 : full_adder port map (N3_9_54,N3_10_54,N3_11_54,N4_6_54,N4_7_55);
-- In matrix 3 adding FA to column 54 
	-- signal N4_8_54 : std_logic;
	-- signal N4_9_55 : std_logic;
	FA1113 : full_adder port map (N3_12_54,N3_13_54,N3_14_54,N4_8_54,N4_9_55);
-- In matrix 3 adding FA to column 54 
	-- signal N4_10_54 : std_logic;
	-- signal N4_11_55 : std_logic;
	FA1114 : full_adder port map (N3_15_54,N3_16_54,N3_17_54,N4_10_54,N4_11_55);
-- In matrix 3 adding FA to column 54 
	-- signal N4_12_54 : std_logic;
	-- signal N4_13_55 : std_logic;
	FA1115 : full_adder port map (N3_18_54,N3_19_54,N3_20_54,N4_12_54,N4_13_55);
-- In matrix 3 adding FA to column 54 
	-- signal N4_14_54 : std_logic;
	-- signal N4_15_55 : std_logic;
	FA1116 : full_adder port map (N3_21_54,N3_22_54,N3_23_54,N4_14_54,N4_15_55);
-- In matrix 3 adding FA to column 55 
	-- signal N4_0_55 : std_logic;
	-- signal N4_1_56 : std_logic;
	FA1117 : full_adder port map (N3_0_55,N3_1_55,N3_2_55,N4_0_55,N4_1_56);
-- In matrix 3 adding FA to column 55 
	-- signal N4_2_55 : std_logic;
	-- signal N4_3_56 : std_logic;
	FA1118 : full_adder port map (N3_3_55,N3_4_55,N3_5_55,N4_2_55,N4_3_56);
-- In matrix 3 adding FA to column 55 
	-- signal N4_4_55 : std_logic;
	-- signal N4_5_56 : std_logic;
	FA1119 : full_adder port map (N3_6_55,N3_7_55,N3_8_55,N4_4_55,N4_5_56);
-- In matrix 3 adding FA to column 55 
	-- signal N4_6_55 : std_logic;
	-- signal N4_7_56 : std_logic;
	FA1120 : full_adder port map (N3_9_55,N3_10_55,N3_11_55,N4_6_55,N4_7_56);
-- In matrix 3 adding FA to column 55 
	-- signal N4_8_55 : std_logic;
	-- signal N4_9_56 : std_logic;
	FA1121 : full_adder port map (N3_12_55,N3_13_55,N3_14_55,N4_8_55,N4_9_56);
-- In matrix 3 adding FA to column 55 
	-- signal N4_10_55 : std_logic;
	-- signal N4_11_56 : std_logic;
	FA1122 : full_adder port map (N3_15_55,N3_16_55,N3_17_55,N4_10_55,N4_11_56);
-- In matrix 3 adding FA to column 55 
	-- signal N4_12_55 : std_logic;
	-- signal N4_13_56 : std_logic;
	FA1123 : full_adder port map (N3_18_55,N3_19_55,N3_20_55,N4_12_55,N4_13_56);
-- In matrix 3 adding FA to column 55 
	-- signal N4_14_55 : std_logic;
	-- signal N4_15_56 : std_logic;
	FA1124 : full_adder port map (N3_21_55,N3_22_55,N3_23_55,N4_14_55,N4_15_56);
-- In matrix 3 adding FA to column 56 
	-- signal N4_0_56 : std_logic;
	-- signal N4_1_57 : std_logic;
	FA1125 : full_adder port map (N3_0_56,N3_1_56,N3_2_56,N4_0_56,N4_1_57);
-- In matrix 3 adding FA to column 56 
	-- signal N4_2_56 : std_logic;
	-- signal N4_3_57 : std_logic;
	FA1126 : full_adder port map (N3_3_56,N3_4_56,N3_5_56,N4_2_56,N4_3_57);
-- In matrix 3 adding FA to column 56 
	-- signal N4_4_56 : std_logic;
	-- signal N4_5_57 : std_logic;
	FA1127 : full_adder port map (N3_6_56,N3_7_56,N3_8_56,N4_4_56,N4_5_57);
-- In matrix 3 adding FA to column 56 
	-- signal N4_6_56 : std_logic;
	-- signal N4_7_57 : std_logic;
	FA1128 : full_adder port map (N3_9_56,N3_10_56,N3_11_56,N4_6_56,N4_7_57);
-- In matrix 3 adding FA to column 56 
	-- signal N4_8_56 : std_logic;
	-- signal N4_9_57 : std_logic;
	FA1129 : full_adder port map (N3_12_56,N3_13_56,N3_14_56,N4_8_56,N4_9_57);
-- In matrix 3 adding FA to column 56 
	-- signal N4_10_56 : std_logic;
	-- signal N4_11_57 : std_logic;
	FA1130 : full_adder port map (N3_15_56,N3_16_56,N3_17_56,N4_10_56,N4_11_57);
-- In matrix 3 adding FA to column 56 
	-- signal N4_12_56 : std_logic;
	-- signal N4_13_57 : std_logic;
	FA1131 : full_adder port map (N3_18_56,N3_19_56,N3_20_56,N4_12_56,N4_13_57);
-- In matrix 3 adding FA to column 56 
	-- signal N4_14_56 : std_logic;
	-- signal N4_15_57 : std_logic;
	FA1132 : full_adder port map (N3_21_56,N3_22_56,N3_23_56,N4_14_56,N4_15_57);
-- In matrix 3 adding FA to column 57 
	-- signal N4_0_57 : std_logic;
	-- signal N4_1_58 : std_logic;
	FA1133 : full_adder port map (N3_0_57,N3_1_57,N3_2_57,N4_0_57,N4_1_58);
-- In matrix 3 adding FA to column 57 
	-- signal N4_2_57 : std_logic;
	-- signal N4_3_58 : std_logic;
	FA1134 : full_adder port map (N3_3_57,N3_4_57,N3_5_57,N4_2_57,N4_3_58);
-- In matrix 3 adding FA to column 57 
	-- signal N4_4_57 : std_logic;
	-- signal N4_5_58 : std_logic;
	FA1135 : full_adder port map (N3_6_57,N3_7_57,N3_8_57,N4_4_57,N4_5_58);
-- In matrix 3 adding FA to column 57 
	-- signal N4_6_57 : std_logic;
	-- signal N4_7_58 : std_logic;
	FA1136 : full_adder port map (N3_9_57,N3_10_57,N3_11_57,N4_6_57,N4_7_58);
-- In matrix 3 adding FA to column 57 
	-- signal N4_8_57 : std_logic;
	-- signal N4_9_58 : std_logic;
	FA1137 : full_adder port map (N3_12_57,N3_13_57,N3_14_57,N4_8_57,N4_9_58);
-- In matrix 3 adding FA to column 57 
	-- signal N4_10_57 : std_logic;
	-- signal N4_11_58 : std_logic;
	FA1138 : full_adder port map (N3_15_57,N3_16_57,N3_17_57,N4_10_57,N4_11_58);
-- In matrix 3 adding FA to column 57 
	-- signal N4_12_57 : std_logic;
	-- signal N4_13_58 : std_logic;
	FA1139 : full_adder port map (N3_18_57,N3_19_57,N3_20_57,N4_12_57,N4_13_58);
-- In matrix 3 adding FA to column 57 
	-- signal N4_14_57 : std_logic;
	-- signal N4_15_58 : std_logic;
	FA1140 : full_adder port map (N3_21_57,N3_22_57,N3_23_57,N4_14_57,N4_15_58);
-- In matrix 3 adding FA to column 58 
	-- signal N4_0_58 : std_logic;
	-- signal N4_1_59 : std_logic;
	FA1141 : full_adder port map (N3_0_58,N3_1_58,N3_2_58,N4_0_58,N4_1_59);
-- In matrix 3 adding FA to column 58 
	-- signal N4_2_58 : std_logic;
	-- signal N4_3_59 : std_logic;
	FA1142 : full_adder port map (N3_3_58,N3_4_58,N3_5_58,N4_2_58,N4_3_59);
-- In matrix 3 adding FA to column 58 
	-- signal N4_4_58 : std_logic;
	-- signal N4_5_59 : std_logic;
	FA1143 : full_adder port map (N3_6_58,N3_7_58,N3_8_58,N4_4_58,N4_5_59);
-- In matrix 3 adding FA to column 58 
	-- signal N4_6_58 : std_logic;
	-- signal N4_7_59 : std_logic;
	FA1144 : full_adder port map (N3_9_58,N3_10_58,N3_11_58,N4_6_58,N4_7_59);
-- In matrix 3 adding FA to column 58 
	-- signal N4_8_58 : std_logic;
	-- signal N4_9_59 : std_logic;
	FA1145 : full_adder port map (N3_12_58,N3_13_58,N3_14_58,N4_8_58,N4_9_59);
-- In matrix 3 adding FA to column 58 
	-- signal N4_10_58 : std_logic;
	-- signal N4_11_59 : std_logic;
	FA1146 : full_adder port map (N3_15_58,N3_16_58,N3_17_58,N4_10_58,N4_11_59);
-- In matrix 3 adding FA to column 58 
	-- signal N4_12_58 : std_logic;
	-- signal N4_13_59 : std_logic;
	FA1147 : full_adder port map (N3_18_58,N3_19_58,N3_20_58,N4_12_58,N4_13_59);
-- In matrix 3 adding FA to column 58 
	-- signal N4_14_58 : std_logic;
	-- signal N4_15_59 : std_logic;
	FA1148 : full_adder port map (N3_21_58,N3_22_58,N3_23_58,N4_14_58,N4_15_59);
-- In matrix 3 adding FA to column 59 
	-- signal N4_0_59 : std_logic;
	-- signal N4_1_60 : std_logic;
	FA1149 : full_adder port map (N3_0_59,N3_1_59,N3_2_59,N4_0_59,N4_1_60);
-- In matrix 3 adding FA to column 59 
	-- signal N4_2_59 : std_logic;
	-- signal N4_3_60 : std_logic;
	FA1150 : full_adder port map (N3_3_59,N3_4_59,N3_5_59,N4_2_59,N4_3_60);
-- In matrix 3 adding FA to column 59 
	-- signal N4_4_59 : std_logic;
	-- signal N4_5_60 : std_logic;
	FA1151 : full_adder port map (N3_6_59,N3_7_59,N3_8_59,N4_4_59,N4_5_60);
-- In matrix 3 adding FA to column 59 
	-- signal N4_6_59 : std_logic;
	-- signal N4_7_60 : std_logic;
	FA1152 : full_adder port map (N3_9_59,N3_10_59,N3_11_59,N4_6_59,N4_7_60);
-- In matrix 3 adding FA to column 59 
	-- signal N4_8_59 : std_logic;
	-- signal N4_9_60 : std_logic;
	FA1153 : full_adder port map (N3_12_59,N3_13_59,N3_14_59,N4_8_59,N4_9_60);
-- In matrix 3 adding FA to column 59 
	-- signal N4_10_59 : std_logic;
	-- signal N4_11_60 : std_logic;
	FA1154 : full_adder port map (N3_15_59,N3_16_59,N3_17_59,N4_10_59,N4_11_60);
-- In matrix 3 adding FA to column 59 
	-- signal N4_12_59 : std_logic;
	-- signal N4_13_60 : std_logic;
	FA1155 : full_adder port map (N3_18_59,N3_19_59,N3_20_59,N4_12_59,N4_13_60);
-- In matrix 3 adding FA to column 59 
	-- signal N4_14_59 : std_logic;
	-- signal N4_15_60 : std_logic;
	FA1156 : full_adder port map (N3_21_59,N3_22_59,N3_23_59,N4_14_59,N4_15_60);
-- In matrix 3 adding FA to column 60 
	-- signal N4_0_60 : std_logic;
	-- signal N4_1_61 : std_logic;
	FA1157 : full_adder port map (N3_0_60,N3_1_60,N3_2_60,N4_0_60,N4_1_61);
-- In matrix 3 adding FA to column 60 
	-- signal N4_2_60 : std_logic;
	-- signal N4_3_61 : std_logic;
	FA1158 : full_adder port map (N3_3_60,N3_4_60,N3_5_60,N4_2_60,N4_3_61);
-- In matrix 3 adding FA to column 60 
	-- signal N4_4_60 : std_logic;
	-- signal N4_5_61 : std_logic;
	FA1159 : full_adder port map (N3_6_60,N3_7_60,N3_8_60,N4_4_60,N4_5_61);
-- In matrix 3 adding FA to column 60 
	-- signal N4_6_60 : std_logic;
	-- signal N4_7_61 : std_logic;
	FA1160 : full_adder port map (N3_9_60,N3_10_60,N3_11_60,N4_6_60,N4_7_61);
-- In matrix 3 adding FA to column 60 
	-- signal N4_8_60 : std_logic;
	-- signal N4_9_61 : std_logic;
	FA1161 : full_adder port map (N3_12_60,N3_13_60,N3_14_60,N4_8_60,N4_9_61);
-- In matrix 3 adding FA to column 60 
	-- signal N4_10_60 : std_logic;
	-- signal N4_11_61 : std_logic;
	FA1162 : full_adder port map (N3_15_60,N3_16_60,N3_17_60,N4_10_60,N4_11_61);
-- In matrix 3 adding FA to column 60 
	-- signal N4_12_60 : std_logic;
	-- signal N4_13_61 : std_logic;
	FA1163 : full_adder port map (N3_18_60,N3_19_60,N3_20_60,N4_12_60,N4_13_61);
-- In matrix 3 adding FA to column 60 
	-- signal N4_14_60 : std_logic;
	-- signal N4_15_61 : std_logic;
	FA1164 : full_adder port map (N3_21_60,N3_22_60,N3_23_60,N4_14_60,N4_15_61);
-- In matrix 3 adding FA to column 61 
	-- signal N4_0_61 : std_logic;
	-- signal N4_1_62 : std_logic;
	FA1165 : full_adder port map (N3_0_61,N3_1_61,N3_2_61,N4_0_61,N4_1_62);
-- In matrix 3 adding FA to column 61 
	-- signal N4_2_61 : std_logic;
	-- signal N4_3_62 : std_logic;
	FA1166 : full_adder port map (N3_3_61,N3_4_61,N3_5_61,N4_2_61,N4_3_62);
-- In matrix 3 adding FA to column 61 
	-- signal N4_4_61 : std_logic;
	-- signal N4_5_62 : std_logic;
	FA1167 : full_adder port map (N3_6_61,N3_7_61,N3_8_61,N4_4_61,N4_5_62);
-- In matrix 3 adding FA to column 61 
	-- signal N4_6_61 : std_logic;
	-- signal N4_7_62 : std_logic;
	FA1168 : full_adder port map (N3_9_61,N3_10_61,N3_11_61,N4_6_61,N4_7_62);
-- In matrix 3 adding FA to column 61 
	-- signal N4_8_61 : std_logic;
	-- signal N4_9_62 : std_logic;
	FA1169 : full_adder port map (N3_12_61,N3_13_61,N3_14_61,N4_8_61,N4_9_62);
-- In matrix 3 adding FA to column 61 
	-- signal N4_10_61 : std_logic;
	-- signal N4_11_62 : std_logic;
	FA1170 : full_adder port map (N3_15_61,N3_16_61,N3_17_61,N4_10_61,N4_11_62);
-- In matrix 3 adding FA to column 61 
	-- signal N4_12_61 : std_logic;
	-- signal N4_13_62 : std_logic;
	FA1171 : full_adder port map (N3_18_61,N3_19_61,N3_20_61,N4_12_61,N4_13_62);
-- In matrix 3 adding FA to column 61 
	-- signal N4_14_61 : std_logic;
	-- signal N4_15_62 : std_logic;
	FA1172 : full_adder port map (N3_21_61,N3_22_61,N3_23_61,N4_14_61,N4_15_62);
-- In matrix 3 adding FA to column 62 
	-- signal N4_0_62 : std_logic;
	-- signal N4_1_63 : std_logic;
	FA1173 : full_adder port map (N3_0_62,N3_1_62,N3_2_62,N4_0_62,N4_1_63);
-- In matrix 3 adding FA to column 62 
	-- signal N4_2_62 : std_logic;
	-- signal N4_3_63 : std_logic;
	FA1174 : full_adder port map (N3_3_62,N3_4_62,N3_5_62,N4_2_62,N4_3_63);
-- In matrix 3 adding FA to column 62 
	-- signal N4_4_62 : std_logic;
	-- signal N4_5_63 : std_logic;
	FA1175 : full_adder port map (N3_6_62,N3_7_62,N3_8_62,N4_4_62,N4_5_63);
-- In matrix 3 adding FA to column 62 
	-- signal N4_6_62 : std_logic;
	-- signal N4_7_63 : std_logic;
	FA1176 : full_adder port map (N3_9_62,N3_10_62,N3_11_62,N4_6_62,N4_7_63);
-- In matrix 3 adding FA to column 62 
	-- signal N4_8_62 : std_logic;
	-- signal N4_9_63 : std_logic;
	FA1177 : full_adder port map (N3_12_62,N3_13_62,N3_14_62,N4_8_62,N4_9_63);
-- In matrix 3 adding FA to column 62 
	-- signal N4_10_62 : std_logic;
	-- signal N4_11_63 : std_logic;
	FA1178 : full_adder port map (N3_15_62,N3_16_62,N3_17_62,N4_10_62,N4_11_63);
-- In matrix 3 adding FA to column 62 
	-- signal N4_12_62 : std_logic;
	-- signal N4_13_63 : std_logic;
	FA1179 : full_adder port map (N3_18_62,N3_19_62,N3_20_62,N4_12_62,N4_13_63);
-- In matrix 3 adding FA to column 62 
	-- signal N4_14_62 : std_logic;
	-- signal N4_15_63 : std_logic;
	FA1180 : full_adder port map (N3_21_62,N3_22_62,N3_23_62,N4_14_62,N4_15_63);
-- In matrix 3 adding FA to column 63 
	-- signal N4_0_63 : std_logic;
	-- signal N4_1_64 : std_logic;
	FA1181 : full_adder port map (N3_0_63,N3_1_63,N3_2_63,N4_0_63,N4_1_64);
-- In matrix 3 adding FA to column 63 
	-- signal N4_2_63 : std_logic;
	-- signal N4_3_64 : std_logic;
	FA1182 : full_adder port map (N3_3_63,N3_4_63,N3_5_63,N4_2_63,N4_3_64);
-- In matrix 3 adding FA to column 63 
	-- signal N4_4_63 : std_logic;
	-- signal N4_5_64 : std_logic;
	FA1183 : full_adder port map (N3_6_63,N3_7_63,N3_8_63,N4_4_63,N4_5_64);
-- In matrix 3 adding FA to column 63 
	-- signal N4_6_63 : std_logic;
	-- signal N4_7_64 : std_logic;
	FA1184 : full_adder port map (N3_9_63,N3_10_63,N3_11_63,N4_6_63,N4_7_64);
-- In matrix 3 adding FA to column 63 
	-- signal N4_8_63 : std_logic;
	-- signal N4_9_64 : std_logic;
	FA1185 : full_adder port map (N3_12_63,N3_13_63,N3_14_63,N4_8_63,N4_9_64);
-- In matrix 3 adding FA to column 63 
	-- signal N4_10_63 : std_logic;
	-- signal N4_11_64 : std_logic;
	FA1186 : full_adder port map (N3_15_63,N3_16_63,N3_17_63,N4_10_63,N4_11_64);
-- In matrix 3 adding FA to column 63 
	-- signal N4_12_63 : std_logic;
	-- signal N4_13_64 : std_logic;
	FA1187 : full_adder port map (N3_18_63,N3_19_63,N3_20_63,N4_12_63,N4_13_64);
-- In matrix 3 adding FA to column 63 
	-- signal N4_14_63 : std_logic;
	-- signal N4_15_64 : std_logic;
	FA1188 : full_adder port map (N3_21_63,N3_22_63,N3_23_63,N4_14_63,N4_15_64);
-- In matrix 3 adding FA to column 64 
	-- signal N4_0_64 : std_logic;
	-- signal N4_1_65 : std_logic;
	FA1189 : full_adder port map (N3_0_64,N3_1_64,N3_2_64,N4_0_64,N4_1_65);
-- In matrix 3 adding FA to column 64 
	-- signal N4_2_64 : std_logic;
	-- signal N4_3_65 : std_logic;
	FA1190 : full_adder port map (N3_3_64,N3_4_64,N3_5_64,N4_2_64,N4_3_65);
-- In matrix 3 adding FA to column 64 
	-- signal N4_4_64 : std_logic;
	-- signal N4_5_65 : std_logic;
	FA1191 : full_adder port map (N3_6_64,N3_7_64,N3_8_64,N4_4_64,N4_5_65);
-- In matrix 3 adding FA to column 64 
	-- signal N4_6_64 : std_logic;
	-- signal N4_7_65 : std_logic;
	FA1192 : full_adder port map (N3_9_64,N3_10_64,N3_11_64,N4_6_64,N4_7_65);
-- In matrix 3 adding FA to column 64 
	-- signal N4_8_64 : std_logic;
	-- signal N4_9_65 : std_logic;
	FA1193 : full_adder port map (N3_12_64,N3_13_64,N3_14_64,N4_8_64,N4_9_65);
-- In matrix 3 adding FA to column 64 
	-- signal N4_10_64 : std_logic;
	-- signal N4_11_65 : std_logic;
	FA1194 : full_adder port map (N3_15_64,N3_16_64,N3_17_64,N4_10_64,N4_11_65);
-- In matrix 3 adding FA to column 64 
	-- signal N4_12_64 : std_logic;
	-- signal N4_13_65 : std_logic;
	FA1195 : full_adder port map (N3_18_64,N3_19_64,N3_20_64,N4_12_64,N4_13_65);
-- In matrix 3 adding FA to column 64 
	-- signal N4_14_64 : std_logic;
	-- signal N4_15_65 : std_logic;
	FA1196 : full_adder port map (N3_21_64,N3_22_64,N3_23_64,N4_14_64,N4_15_65);
-- In matrix 3 adding FA to column 65 
	-- signal N4_0_65 : std_logic;
	-- signal N4_1_66 : std_logic;
	FA1197 : full_adder port map (N3_0_65,N3_1_65,N3_2_65,N4_0_65,N4_1_66);
-- In matrix 3 adding FA to column 65 
	-- signal N4_2_65 : std_logic;
	-- signal N4_3_66 : std_logic;
	FA1198 : full_adder port map (N3_3_65,N3_4_65,N3_5_65,N4_2_65,N4_3_66);
-- In matrix 3 adding FA to column 65 
	-- signal N4_4_65 : std_logic;
	-- signal N4_5_66 : std_logic;
	FA1199 : full_adder port map (N3_6_65,N3_7_65,N3_8_65,N4_4_65,N4_5_66);
-- In matrix 3 adding FA to column 65 
	-- signal N4_6_65 : std_logic;
	-- signal N4_7_66 : std_logic;
	FA1200 : full_adder port map (N3_9_65,N3_10_65,N3_11_65,N4_6_65,N4_7_66);
-- In matrix 3 adding FA to column 65 
	-- signal N4_8_65 : std_logic;
	-- signal N4_9_66 : std_logic;
	FA1201 : full_adder port map (N3_12_65,N3_13_65,N3_14_65,N4_8_65,N4_9_66);
-- In matrix 3 adding FA to column 65 
	-- signal N4_10_65 : std_logic;
	-- signal N4_11_66 : std_logic;
	FA1202 : full_adder port map (N3_15_65,N3_16_65,N3_17_65,N4_10_65,N4_11_66);
-- In matrix 3 adding FA to column 65 
	-- signal N4_12_65 : std_logic;
	-- signal N4_13_66 : std_logic;
	FA1203 : full_adder port map (N3_18_65,N3_19_65,N3_20_65,N4_12_65,N4_13_66);
-- In matrix 3 adding FA to column 65 
	-- signal N4_14_65 : std_logic;
	-- signal N4_15_66 : std_logic;
	FA1204 : full_adder port map (N3_21_65,N3_22_65,N3_23_65,N4_14_65,N4_15_66);
-- In matrix 3 adding FA to column 66 
	-- signal N4_0_66 : std_logic;
	-- signal N4_1_67 : std_logic;
	FA1205 : full_adder port map (N3_0_66,N3_1_66,N3_2_66,N4_0_66,N4_1_67);
-- In matrix 3 adding FA to column 66 
	-- signal N4_2_66 : std_logic;
	-- signal N4_3_67 : std_logic;
	FA1206 : full_adder port map (N3_3_66,N3_4_66,N3_5_66,N4_2_66,N4_3_67);
-- In matrix 3 adding FA to column 66 
	-- signal N4_4_66 : std_logic;
	-- signal N4_5_67 : std_logic;
	FA1207 : full_adder port map (N3_6_66,N3_7_66,N3_8_66,N4_4_66,N4_5_67);
-- In matrix 3 adding FA to column 66 
	-- signal N4_6_66 : std_logic;
	-- signal N4_7_67 : std_logic;
	FA1208 : full_adder port map (N3_9_66,N3_10_66,N3_11_66,N4_6_66,N4_7_67);
-- In matrix 3 adding FA to column 66 
	-- signal N4_8_66 : std_logic;
	-- signal N4_9_67 : std_logic;
	FA1209 : full_adder port map (N3_12_66,N3_13_66,N3_14_66,N4_8_66,N4_9_67);
-- In matrix 3 adding FA to column 66 
	-- signal N4_10_66 : std_logic;
	-- signal N4_11_67 : std_logic;
	FA1210 : full_adder port map (N3_15_66,N3_16_66,N3_17_66,N4_10_66,N4_11_67);
-- In matrix 3 adding FA to column 66 
	-- signal N4_12_66 : std_logic;
	-- signal N4_13_67 : std_logic;
	FA1211 : full_adder port map (N3_18_66,N3_19_66,N3_20_66,N4_12_66,N4_13_67);
-- In matrix 3 adding FA to column 66 
	-- signal N4_14_66 : std_logic;
	-- signal N4_15_67 : std_logic;
	FA1212 : full_adder port map (N3_21_66,N3_22_66,N3_23_66,N4_14_66,N4_15_67);
-- In matrix 3 adding FA to column 67 
	-- signal N4_0_67 : std_logic;
	-- signal N4_1_68 : std_logic;
	FA1213 : full_adder port map (N3_0_67,N3_1_67,N3_2_67,N4_0_67,N4_1_68);
-- In matrix 3 adding FA to column 67 
	-- signal N4_2_67 : std_logic;
	-- signal N4_3_68 : std_logic;
	FA1214 : full_adder port map (N3_3_67,N3_4_67,N3_5_67,N4_2_67,N4_3_68);
-- In matrix 3 adding FA to column 67 
	-- signal N4_4_67 : std_logic;
	-- signal N4_5_68 : std_logic;
	FA1215 : full_adder port map (N3_6_67,N3_7_67,N3_8_67,N4_4_67,N4_5_68);
-- In matrix 3 adding FA to column 67 
	-- signal N4_6_67 : std_logic;
	-- signal N4_7_68 : std_logic;
	FA1216 : full_adder port map (N3_9_67,N3_10_67,N3_11_67,N4_6_67,N4_7_68);
-- In matrix 3 adding FA to column 67 
	-- signal N4_8_67 : std_logic;
	-- signal N4_9_68 : std_logic;
	FA1217 : full_adder port map (N3_12_67,N3_13_67,N3_14_67,N4_8_67,N4_9_68);
-- In matrix 3 adding FA to column 67 
	-- signal N4_10_67 : std_logic;
	-- signal N4_11_68 : std_logic;
	FA1218 : full_adder port map (N3_15_67,N3_16_67,N3_17_67,N4_10_67,N4_11_68);
-- In matrix 3 adding FA to column 67 
	-- signal N4_12_67 : std_logic;
	-- signal N4_13_68 : std_logic;
	FA1219 : full_adder port map (N3_18_67,N3_19_67,N3_20_67,N4_12_67,N4_13_68);
-- In matrix 3 adding FA to column 67 
	-- signal N4_14_67 : std_logic;
	-- signal N4_15_68 : std_logic;
	FA1220 : full_adder port map (N3_21_67,N3_22_67,N3_23_67,N4_14_67,N4_15_68);
-- In matrix 3 adding FA to column 68 
	-- signal N4_0_68 : std_logic;
	-- signal N4_1_69 : std_logic;
	FA1221 : full_adder port map (N3_0_68,N3_1_68,N3_2_68,N4_0_68,N4_1_69);
-- In matrix 3 adding FA to column 68 
	-- signal N4_2_68 : std_logic;
	-- signal N4_3_69 : std_logic;
	FA1222 : full_adder port map (N3_3_68,N3_4_68,N3_5_68,N4_2_68,N4_3_69);
-- In matrix 3 adding FA to column 68 
	-- signal N4_4_68 : std_logic;
	-- signal N4_5_69 : std_logic;
	FA1223 : full_adder port map (N3_6_68,N3_7_68,N3_8_68,N4_4_68,N4_5_69);
-- In matrix 3 adding FA to column 68 
	-- signal N4_6_68 : std_logic;
	-- signal N4_7_69 : std_logic;
	FA1224 : full_adder port map (N3_9_68,N3_10_68,N3_11_68,N4_6_68,N4_7_69);
-- In matrix 3 adding FA to column 68 
	-- signal N4_8_68 : std_logic;
	-- signal N4_9_69 : std_logic;
	FA1225 : full_adder port map (N3_12_68,N3_13_68,N3_14_68,N4_8_68,N4_9_69);
-- In matrix 3 adding FA to column 68 
	-- signal N4_10_68 : std_logic;
	-- signal N4_11_69 : std_logic;
	FA1226 : full_adder port map (N3_15_68,N3_16_68,N3_17_68,N4_10_68,N4_11_69);
-- In matrix 3 adding FA to column 68 
	-- signal N4_12_68 : std_logic;
	-- signal N4_13_69 : std_logic;
	FA1227 : full_adder port map (N3_18_68,N3_19_68,N3_20_68,N4_12_68,N4_13_69);
-- In matrix 3 adding FA to column 68 
	-- signal N4_14_68 : std_logic;
	-- signal N4_15_69 : std_logic;
	FA1228 : full_adder port map (N3_21_68,N3_22_68,N3_23_68,N4_14_68,N4_15_69);
-- In matrix 3 adding FA to column 69 
	-- signal N4_0_69 : std_logic;
	-- signal N4_1_70 : std_logic;
	FA1229 : full_adder port map (N3_0_69,N3_1_69,N3_2_69,N4_0_69,N4_1_70);
-- In matrix 3 adding FA to column 69 
	-- signal N4_2_69 : std_logic;
	-- signal N4_3_70 : std_logic;
	FA1230 : full_adder port map (N3_3_69,N3_4_69,N3_5_69,N4_2_69,N4_3_70);
-- In matrix 3 adding FA to column 69 
	-- signal N4_4_69 : std_logic;
	-- signal N4_5_70 : std_logic;
	FA1231 : full_adder port map (N3_6_69,N3_7_69,N3_8_69,N4_4_69,N4_5_70);
-- In matrix 3 adding FA to column 69 
	-- signal N4_6_69 : std_logic;
	-- signal N4_7_70 : std_logic;
	FA1232 : full_adder port map (N3_9_69,N3_10_69,N3_11_69,N4_6_69,N4_7_70);
-- In matrix 3 adding FA to column 69 
	-- signal N4_8_69 : std_logic;
	-- signal N4_9_70 : std_logic;
	FA1233 : full_adder port map (N3_12_69,N3_13_69,N3_14_69,N4_8_69,N4_9_70);
-- In matrix 3 adding FA to column 69 
	-- signal N4_10_69 : std_logic;
	-- signal N4_11_70 : std_logic;
	FA1234 : full_adder port map (N3_15_69,N3_16_69,N3_17_69,N4_10_69,N4_11_70);
-- In matrix 3 adding FA to column 69 
	-- signal N4_12_69 : std_logic;
	-- signal N4_13_70 : std_logic;
	FA1235 : full_adder port map (N3_18_69,N3_19_69,N3_20_69,N4_12_69,N4_13_70);
-- In matrix 3 adding FA to column 69 
	-- signal N4_14_69 : std_logic;
	-- signal N4_15_70 : std_logic;
	FA1236 : full_adder port map (N3_21_69,N3_22_69,N3_23_69,N4_14_69,N4_15_70);
-- In matrix 3 adding FA to column 70 
	-- signal N4_0_70 : std_logic;
	-- signal N4_1_71 : std_logic;
	FA1237 : full_adder port map (N3_0_70,N3_1_70,N3_2_70,N4_0_70,N4_1_71);
-- In matrix 3 adding FA to column 70 
	-- signal N4_2_70 : std_logic;
	-- signal N4_3_71 : std_logic;
	FA1238 : full_adder port map (N3_3_70,N3_4_70,N3_5_70,N4_2_70,N4_3_71);
-- In matrix 3 adding FA to column 70 
	-- signal N4_4_70 : std_logic;
	-- signal N4_5_71 : std_logic;
	FA1239 : full_adder port map (N3_6_70,N3_7_70,N3_8_70,N4_4_70,N4_5_71);
-- In matrix 3 adding FA to column 70 
	-- signal N4_6_70 : std_logic;
	-- signal N4_7_71 : std_logic;
	FA1240 : full_adder port map (N3_9_70,N3_10_70,N3_11_70,N4_6_70,N4_7_71);
-- In matrix 3 adding FA to column 70 
	-- signal N4_8_70 : std_logic;
	-- signal N4_9_71 : std_logic;
	FA1241 : full_adder port map (N3_12_70,N3_13_70,N3_14_70,N4_8_70,N4_9_71);
-- In matrix 3 adding FA to column 70 
	-- signal N4_10_70 : std_logic;
	-- signal N4_11_71 : std_logic;
	FA1242 : full_adder port map (N3_15_70,N3_16_70,N3_17_70,N4_10_70,N4_11_71);
-- In matrix 3 adding FA to column 70 
	-- signal N4_12_70 : std_logic;
	-- signal N4_13_71 : std_logic;
	FA1243 : full_adder port map (N3_18_70,N3_19_70,N3_20_70,N4_12_70,N4_13_71);
-- In matrix 3 adding FA to column 70 
	-- signal N4_14_70 : std_logic;
	-- signal N4_15_71 : std_logic;
	FA1244 : full_adder port map (N3_21_70,N3_22_70,N3_23_70,N4_14_70,N4_15_71);
-- In matrix 3 adding FA to column 71 
	-- signal N4_0_71 : std_logic;
	-- signal N4_1_72 : std_logic;
	FA1245 : full_adder port map (N0_52_71,N3_0_71,N3_1_71,N4_0_71,N4_1_72);
-- In matrix 3 adding FA to column 71 
	-- signal N4_2_71 : std_logic;
	-- signal N4_3_72 : std_logic;
	FA1246 : full_adder port map (N3_2_71,N3_3_71,N3_4_71,N4_2_71,N4_3_72);
-- In matrix 3 adding FA to column 71 
	-- signal N4_4_71 : std_logic;
	-- signal N4_5_72 : std_logic;
	FA1247 : full_adder port map (N3_5_71,N3_6_71,N3_7_71,N4_4_71,N4_5_72);
-- In matrix 3 adding FA to column 71 
	-- signal N4_6_71 : std_logic;
	-- signal N4_7_72 : std_logic;
	FA1248 : full_adder port map (N3_8_71,N3_9_71,N3_10_71,N4_6_71,N4_7_72);
-- In matrix 3 adding FA to column 71 
	-- signal N4_8_71 : std_logic;
	-- signal N4_9_72 : std_logic;
	FA1249 : full_adder port map (N3_11_71,N3_12_71,N3_13_71,N4_8_71,N4_9_72);
-- In matrix 3 adding FA to column 71 
	-- signal N4_10_71 : std_logic;
	-- signal N4_11_72 : std_logic;
	FA1250 : full_adder port map (N3_14_71,N3_15_71,N3_16_71,N4_10_71,N4_11_72);
-- In matrix 3 adding FA to column 71 
	-- signal N4_12_71 : std_logic;
	-- signal N4_13_72 : std_logic;
	FA1251 : full_adder port map (N3_17_71,N3_18_71,N3_19_71,N4_12_71,N4_13_72);
-- In matrix 3 adding FA to column 71 
	-- signal N4_14_71 : std_logic;
	-- signal N4_15_72 : std_logic;
	FA1252 : full_adder port map (N3_20_71,N3_21_71,N3_23_71,N4_14_71,N4_15_72);
-- In matrix 3 adding FA to column 72 
	-- signal N4_0_72 : std_logic;
	-- signal N4_1_73 : std_logic;
	FA1253 : full_adder port map (N0_50_72,N0_51_72,N0_52_72,N4_0_72,N4_1_73);
-- In matrix 3 adding FA to column 72 
	-- signal N4_2_72 : std_logic;
	-- signal N4_3_73 : std_logic;
	FA1254 : full_adder port map (N3_0_72,N3_1_72,N3_2_72,N4_2_72,N4_3_73);
-- In matrix 3 adding FA to column 72 
	-- signal N4_4_72 : std_logic;
	-- signal N4_5_73 : std_logic;
	FA1255 : full_adder port map (N3_3_72,N3_4_72,N3_5_72,N4_4_72,N4_5_73);
-- In matrix 3 adding FA to column 72 
	-- signal N4_6_72 : std_logic;
	-- signal N4_7_73 : std_logic;
	FA1256 : full_adder port map (N3_6_72,N3_7_72,N3_8_72,N4_6_72,N4_7_73);
-- In matrix 3 adding FA to column 72 
	-- signal N4_8_72 : std_logic;
	-- signal N4_9_73 : std_logic;
	FA1257 : full_adder port map (N3_9_72,N3_10_72,N3_11_72,N4_8_72,N4_9_73);
-- In matrix 3 adding FA to column 72 
	-- signal N4_10_72 : std_logic;
	-- signal N4_11_73 : std_logic;
	FA1258 : full_adder port map (N3_12_72,N3_13_72,N3_14_72,N4_10_72,N4_11_73);
-- In matrix 3 adding FA to column 72 
	-- signal N4_12_72 : std_logic;
	-- signal N4_13_73 : std_logic;
	FA1259 : full_adder port map (N3_15_72,N3_16_72,N3_17_72,N4_12_72,N4_13_73);
-- In matrix 3 adding FA to column 72 
	-- signal N4_14_72 : std_logic;
	-- signal N4_15_73 : std_logic;
	FA1260 : full_adder port map (N3_18_72,N3_19_72,N3_21_72,N4_14_72,N4_15_73);
-- In matrix 3 adding FA to column 73 
	-- signal N4_0_73 : std_logic;
	-- signal N4_1_74 : std_logic;
	FA1261 : full_adder port map (N0_48_73,N0_49_73,N0_50_73,N4_0_73,N4_1_74);
-- In matrix 3 adding FA to column 73 
	-- signal N4_2_73 : std_logic;
	-- signal N4_3_74 : std_logic;
	FA1262 : full_adder port map (N0_51_73,N0_52_73,N3_0_73,N4_2_73,N4_3_74);
-- In matrix 3 adding FA to column 73 
	-- signal N4_4_73 : std_logic;
	-- signal N4_5_74 : std_logic;
	FA1263 : full_adder port map (N3_1_73,N3_2_73,N3_3_73,N4_4_73,N4_5_74);
-- In matrix 3 adding FA to column 73 
	-- signal N4_6_73 : std_logic;
	-- signal N4_7_74 : std_logic;
	FA1264 : full_adder port map (N3_4_73,N3_5_73,N3_6_73,N4_6_73,N4_7_74);
-- In matrix 3 adding FA to column 73 
	-- signal N4_8_73 : std_logic;
	-- signal N4_9_74 : std_logic;
	FA1265 : full_adder port map (N3_7_73,N3_8_73,N3_9_73,N4_8_73,N4_9_74);
-- In matrix 3 adding FA to column 73 
	-- signal N4_10_73 : std_logic;
	-- signal N4_11_74 : std_logic;
	FA1266 : full_adder port map (N3_10_73,N3_11_73,N3_12_73,N4_10_73,N4_11_74);
-- In matrix 3 adding FA to column 73 
	-- signal N4_12_73 : std_logic;
	-- signal N4_13_74 : std_logic;
	FA1267 : full_adder port map (N3_13_73,N3_14_73,N3_15_73,N4_12_73,N4_13_74);
-- In matrix 3 adding FA to column 73 
	-- signal N4_14_73 : std_logic;
	-- signal N4_15_74 : std_logic;
	FA1268 : full_adder port map (N3_16_73,N3_17_73,N3_19_73,N4_14_73,N4_15_74);
-- In matrix 3 adding FA to column 74 
	-- signal N4_0_74 : std_logic;
	-- signal N4_1_75 : std_logic;
	FA1269 : full_adder port map (N0_46_74,N0_47_74,N0_48_74,N4_0_74,N4_1_75);
-- In matrix 3 adding FA to column 74 
	-- signal N4_2_74 : std_logic;
	-- signal N4_3_75 : std_logic;
	FA1270 : full_adder port map (N0_49_74,N0_50_74,N0_51_74,N4_2_74,N4_3_75);
-- In matrix 3 adding FA to column 74 
	-- signal N4_4_74 : std_logic;
	-- signal N4_5_75 : std_logic;
	FA1271 : full_adder port map (N0_52_74,N3_0_74,N3_1_74,N4_4_74,N4_5_75);
-- In matrix 3 adding FA to column 74 
	-- signal N4_6_74 : std_logic;
	-- signal N4_7_75 : std_logic;
	FA1272 : full_adder port map (N3_2_74,N3_3_74,N3_4_74,N4_6_74,N4_7_75);
-- In matrix 3 adding FA to column 74 
	-- signal N4_8_74 : std_logic;
	-- signal N4_9_75 : std_logic;
	FA1273 : full_adder port map (N3_5_74,N3_6_74,N3_7_74,N4_8_74,N4_9_75);
-- In matrix 3 adding FA to column 74 
	-- signal N4_10_74 : std_logic;
	-- signal N4_11_75 : std_logic;
	FA1274 : full_adder port map (N3_8_74,N3_9_74,N3_10_74,N4_10_74,N4_11_75);
-- In matrix 3 adding FA to column 74 
	-- signal N4_12_74 : std_logic;
	-- signal N4_13_75 : std_logic;
	FA1275 : full_adder port map (N3_11_74,N3_12_74,N3_13_74,N4_12_74,N4_13_75);
-- In matrix 3 adding FA to column 74 
	-- signal N4_14_74 : std_logic;
	-- signal N4_15_75 : std_logic;
	FA1276 : full_adder port map (N3_14_74,N3_15_74,N3_17_74,N4_14_74,N4_15_75);
-- In matrix 3 adding FA to column 75 
	-- signal N4_0_75 : std_logic;
	-- signal N4_1_76 : std_logic;
	FA1277 : full_adder port map (N0_44_75,N0_45_75,N0_46_75,N4_0_75,N4_1_76);
-- In matrix 3 adding FA to column 75 
	-- signal N4_2_75 : std_logic;
	-- signal N4_3_76 : std_logic;
	FA1278 : full_adder port map (N0_47_75,N0_48_75,N0_49_75,N4_2_75,N4_3_76);
-- In matrix 3 adding FA to column 75 
	-- signal N4_4_75 : std_logic;
	-- signal N4_5_76 : std_logic;
	FA1279 : full_adder port map (N0_50_75,N0_51_75,N0_52_75,N4_4_75,N4_5_76);
-- In matrix 3 adding FA to column 75 
	-- signal N4_6_75 : std_logic;
	-- signal N4_7_76 : std_logic;
	FA1280 : full_adder port map (N3_0_75,N3_1_75,N3_2_75,N4_6_75,N4_7_76);
-- In matrix 3 adding FA to column 75 
	-- signal N4_8_75 : std_logic;
	-- signal N4_9_76 : std_logic;
	FA1281 : full_adder port map (N3_3_75,N3_4_75,N3_5_75,N4_8_75,N4_9_76);
-- In matrix 3 adding FA to column 75 
	-- signal N4_10_75 : std_logic;
	-- signal N4_11_76 : std_logic;
	FA1282 : full_adder port map (N3_6_75,N3_7_75,N3_8_75,N4_10_75,N4_11_76);
-- In matrix 3 adding FA to column 75 
	-- signal N4_12_75 : std_logic;
	-- signal N4_13_76 : std_logic;
	FA1283 : full_adder port map (N3_9_75,N3_10_75,N3_11_75,N4_12_75,N4_13_76);
-- In matrix 3 adding FA to column 75 
	-- signal N4_14_75 : std_logic;
	-- signal N4_15_76 : std_logic;
	FA1284 : full_adder port map (N3_12_75,N3_13_75,N3_15_75,N4_14_75,N4_15_76);
-- In matrix 3 adding FA to column 76 
	-- signal N4_0_76 : std_logic;
	-- signal N4_1_77 : std_logic;
	FA1285 : full_adder port map (N0_42_76,N0_43_76,N0_44_76,N4_0_76,N4_1_77);
-- In matrix 3 adding FA to column 76 
	-- signal N4_2_76 : std_logic;
	-- signal N4_3_77 : std_logic;
	FA1286 : full_adder port map (N0_45_76,N0_46_76,N0_47_76,N4_2_76,N4_3_77);
-- In matrix 3 adding FA to column 76 
	-- signal N4_4_76 : std_logic;
	-- signal N4_5_77 : std_logic;
	FA1287 : full_adder port map (N0_48_76,N0_49_76,N0_50_76,N4_4_76,N4_5_77);
-- In matrix 3 adding FA to column 76 
	-- signal N4_6_76 : std_logic;
	-- signal N4_7_77 : std_logic;
	FA1288 : full_adder port map (N0_51_76,N0_52_76,N3_0_76,N4_6_76,N4_7_77);
-- In matrix 3 adding FA to column 76 
	-- signal N4_8_76 : std_logic;
	-- signal N4_9_77 : std_logic;
	FA1289 : full_adder port map (N3_1_76,N3_2_76,N3_3_76,N4_8_76,N4_9_77);
-- In matrix 3 adding FA to column 76 
	-- signal N4_10_76 : std_logic;
	-- signal N4_11_77 : std_logic;
	FA1290 : full_adder port map (N3_4_76,N3_5_76,N3_6_76,N4_10_76,N4_11_77);
-- In matrix 3 adding FA to column 76 
	-- signal N4_12_76 : std_logic;
	-- signal N4_13_77 : std_logic;
	FA1291 : full_adder port map (N3_7_76,N3_8_76,N3_9_76,N4_12_76,N4_13_77);
-- In matrix 3 adding FA to column 76 
	-- signal N4_14_76 : std_logic;
	-- signal N4_15_77 : std_logic;
	FA1292 : full_adder port map (N3_10_76,N3_11_76,N3_13_76,N4_14_76,N4_15_77);
-- In matrix 3 adding FA to column 77 
	-- signal N4_0_77 : std_logic;
	-- signal N4_1_78 : std_logic;
	FA1293 : full_adder port map (N0_40_77,N0_41_77,N0_42_77,N4_0_77,N4_1_78);
-- In matrix 3 adding FA to column 77 
	-- signal N4_2_77 : std_logic;
	-- signal N4_3_78 : std_logic;
	FA1294 : full_adder port map (N0_43_77,N0_44_77,N0_45_77,N4_2_77,N4_3_78);
-- In matrix 3 adding FA to column 77 
	-- signal N4_4_77 : std_logic;
	-- signal N4_5_78 : std_logic;
	FA1295 : full_adder port map (N0_46_77,N0_47_77,N0_48_77,N4_4_77,N4_5_78);
-- In matrix 3 adding FA to column 77 
	-- signal N4_6_77 : std_logic;
	-- signal N4_7_78 : std_logic;
	FA1296 : full_adder port map (N0_49_77,N0_50_77,N0_51_77,N4_6_77,N4_7_78);
-- In matrix 3 adding FA to column 77 
	-- signal N4_8_77 : std_logic;
	-- signal N4_9_78 : std_logic;
	FA1297 : full_adder port map (N0_52_77,N3_0_77,N3_1_77,N4_8_77,N4_9_78);
-- In matrix 3 adding FA to column 77 
	-- signal N4_10_77 : std_logic;
	-- signal N4_11_78 : std_logic;
	FA1298 : full_adder port map (N3_2_77,N3_3_77,N3_4_77,N4_10_77,N4_11_78);
-- In matrix 3 adding FA to column 77 
	-- signal N4_12_77 : std_logic;
	-- signal N4_13_78 : std_logic;
	FA1299 : full_adder port map (N3_5_77,N3_6_77,N3_7_77,N4_12_77,N4_13_78);
-- In matrix 3 adding FA to column 77 
	-- signal N4_14_77 : std_logic;
	-- signal N4_15_78 : std_logic;
	FA1300 : full_adder port map (N3_8_77,N3_9_77,N3_11_77,N4_14_77,N4_15_78);
-- In matrix 3 adding FA to column 78 
	-- signal N4_0_78 : std_logic;
	-- signal N4_1_79 : std_logic;
	FA1301 : full_adder port map (N0_38_78,N0_39_78,N0_40_78,N4_0_78,N4_1_79);
-- In matrix 3 adding FA to column 78 
	-- signal N4_2_78 : std_logic;
	-- signal N4_3_79 : std_logic;
	FA1302 : full_adder port map (N0_41_78,N0_42_78,N0_43_78,N4_2_78,N4_3_79);
-- In matrix 3 adding FA to column 78 
	-- signal N4_4_78 : std_logic;
	-- signal N4_5_79 : std_logic;
	FA1303 : full_adder port map (N0_44_78,N0_45_78,N0_46_78,N4_4_78,N4_5_79);
-- In matrix 3 adding FA to column 78 
	-- signal N4_6_78 : std_logic;
	-- signal N4_7_79 : std_logic;
	FA1304 : full_adder port map (N0_47_78,N0_48_78,N0_49_78,N4_6_78,N4_7_79);
-- In matrix 3 adding FA to column 78 
	-- signal N4_8_78 : std_logic;
	-- signal N4_9_79 : std_logic;
	FA1305 : full_adder port map (N0_50_78,N0_51_78,N0_52_78,N4_8_78,N4_9_79);
-- In matrix 3 adding FA to column 78 
	-- signal N4_10_78 : std_logic;
	-- signal N4_11_79 : std_logic;
	FA1306 : full_adder port map (N3_0_78,N3_1_78,N3_2_78,N4_10_78,N4_11_79);
-- In matrix 3 adding FA to column 78 
	-- signal N4_12_78 : std_logic;
	-- signal N4_13_79 : std_logic;
	FA1307 : full_adder port map (N3_3_78,N3_4_78,N3_5_78,N4_12_78,N4_13_79);
-- In matrix 3 adding FA to column 78 
	-- signal N4_14_78 : std_logic;
	-- signal N4_15_79 : std_logic;
	FA1308 : full_adder port map (N3_6_78,N3_7_78,N3_9_78,N4_14_78,N4_15_79);
-- In matrix 3 adding FA to column 79 
	-- signal N4_0_79 : std_logic;
	-- signal N4_1_80 : std_logic;
	FA1309 : full_adder port map (N0_36_79,N0_37_79,N0_38_79,N4_0_79,N4_1_80);
-- In matrix 3 adding FA to column 79 
	-- signal N4_2_79 : std_logic;
	-- signal N4_3_80 : std_logic;
	FA1310 : full_adder port map (N0_39_79,N0_40_79,N0_41_79,N4_2_79,N4_3_80);
-- In matrix 3 adding FA to column 79 
	-- signal N4_4_79 : std_logic;
	-- signal N4_5_80 : std_logic;
	FA1311 : full_adder port map (N0_42_79,N0_43_79,N0_44_79,N4_4_79,N4_5_80);
-- In matrix 3 adding FA to column 79 
	-- signal N4_6_79 : std_logic;
	-- signal N4_7_80 : std_logic;
	FA1312 : full_adder port map (N0_45_79,N0_46_79,N0_47_79,N4_6_79,N4_7_80);
-- In matrix 3 adding FA to column 79 
	-- signal N4_8_79 : std_logic;
	-- signal N4_9_80 : std_logic;
	FA1313 : full_adder port map (N0_48_79,N0_49_79,N0_50_79,N4_8_79,N4_9_80);
-- In matrix 3 adding FA to column 79 
	-- signal N4_10_79 : std_logic;
	-- signal N4_11_80 : std_logic;
	FA1314 : full_adder port map (N0_51_79,N0_52_79,N3_0_79,N4_10_79,N4_11_80);
-- In matrix 3 adding FA to column 79 
	-- signal N4_12_79 : std_logic;
	-- signal N4_13_80 : std_logic;
	FA1315 : full_adder port map (N3_1_79,N3_2_79,N3_3_79,N4_12_79,N4_13_80);
-- In matrix 3 adding FA to column 79 
	-- signal N4_14_79 : std_logic;
	-- signal N4_15_80 : std_logic;
	FA1316 : full_adder port map (N3_4_79,N3_5_79,N3_7_79,N4_14_79,N4_15_80);
-- In matrix 3 adding FA to column 80 
	-- signal N4_0_80 : std_logic;
	-- signal N4_1_81 : std_logic;
	FA1317 : full_adder port map (N0_34_80,N0_35_80,N0_36_80,N4_0_80,N4_1_81);
-- In matrix 3 adding FA to column 80 
	-- signal N4_2_80 : std_logic;
	-- signal N4_3_81 : std_logic;
	FA1318 : full_adder port map (N0_37_80,N0_38_80,N0_39_80,N4_2_80,N4_3_81);
-- In matrix 3 adding FA to column 80 
	-- signal N4_4_80 : std_logic;
	-- signal N4_5_81 : std_logic;
	FA1319 : full_adder port map (N0_40_80,N0_41_80,N0_42_80,N4_4_80,N4_5_81);
-- In matrix 3 adding FA to column 80 
	-- signal N4_6_80 : std_logic;
	-- signal N4_7_81 : std_logic;
	FA1320 : full_adder port map (N0_43_80,N0_44_80,N0_45_80,N4_6_80,N4_7_81);
-- In matrix 3 adding FA to column 80 
	-- signal N4_8_80 : std_logic;
	-- signal N4_9_81 : std_logic;
	FA1321 : full_adder port map (N0_46_80,N0_47_80,N0_48_80,N4_8_80,N4_9_81);
-- In matrix 3 adding FA to column 80 
	-- signal N4_10_80 : std_logic;
	-- signal N4_11_81 : std_logic;
	FA1322 : full_adder port map (N0_49_80,N0_50_80,N0_51_80,N4_10_80,N4_11_81);
-- In matrix 3 adding FA to column 80 
	-- signal N4_12_80 : std_logic;
	-- signal N4_13_81 : std_logic;
	FA1323 : full_adder port map (N0_52_80,N3_0_80,N3_1_80,N4_12_80,N4_13_81);
-- In matrix 3 adding FA to column 80 
	-- signal N4_14_80 : std_logic;
	-- signal N4_15_81 : std_logic;
	FA1324 : full_adder port map (N3_2_80,N3_3_80,N3_5_80,N4_14_80,N4_15_81);
-- In matrix 3 adding FA to column 81 
	-- signal N4_0_81 : std_logic;
	-- signal N4_1_82 : std_logic;
	FA1325 : full_adder port map (N0_32_81,N0_33_81,N0_34_81,N4_0_81,N4_1_82);
-- In matrix 3 adding FA to column 81 
	-- signal N4_2_81 : std_logic;
	-- signal N4_3_82 : std_logic;
	FA1326 : full_adder port map (N0_35_81,N0_36_81,N0_37_81,N4_2_81,N4_3_82);
-- In matrix 3 adding FA to column 81 
	-- signal N4_4_81 : std_logic;
	-- signal N4_5_82 : std_logic;
	FA1327 : full_adder port map (N0_38_81,N0_39_81,N0_40_81,N4_4_81,N4_5_82);
-- In matrix 3 adding FA to column 81 
	-- signal N4_6_81 : std_logic;
	-- signal N4_7_82 : std_logic;
	FA1328 : full_adder port map (N0_41_81,N0_42_81,N0_43_81,N4_6_81,N4_7_82);
-- In matrix 3 adding FA to column 81 
	-- signal N4_8_81 : std_logic;
	-- signal N4_9_82 : std_logic;
	FA1329 : full_adder port map (N0_44_81,N0_45_81,N0_46_81,N4_8_81,N4_9_82);
-- In matrix 3 adding FA to column 81 
	-- signal N4_10_81 : std_logic;
	-- signal N4_11_82 : std_logic;
	FA1330 : full_adder port map (N0_47_81,N0_48_81,N0_49_81,N4_10_81,N4_11_82);
-- In matrix 3 adding FA to column 81 
	-- signal N4_12_81 : std_logic;
	-- signal N4_13_82 : std_logic;
	FA1331 : full_adder port map (N0_50_81,N0_51_81,N0_52_81,N4_12_81,N4_13_82);
-- In matrix 3 adding FA to column 81 
	-- signal N4_14_81 : std_logic;
	-- signal N4_15_82 : std_logic;
	FA1332 : full_adder port map (N3_0_81,N3_1_81,N3_3_81,N4_14_81,N4_15_82);
-- In matrix 3 adding FA to column 82 
	-- signal N4_0_82 : std_logic;
	-- signal N4_1_83 : std_logic;
	FA1333 : full_adder port map (N0_30_82,N0_31_82,N0_32_82,N4_0_82,N4_1_83);
-- In matrix 3 adding FA to column 82 
	-- signal N4_2_82 : std_logic;
	-- signal N4_3_83 : std_logic;
	FA1334 : full_adder port map (N0_33_82,N0_34_82,N0_35_82,N4_2_82,N4_3_83);
-- In matrix 3 adding FA to column 82 
	-- signal N4_4_82 : std_logic;
	-- signal N4_5_83 : std_logic;
	FA1335 : full_adder port map (N0_36_82,N0_37_82,N0_38_82,N4_4_82,N4_5_83);
-- In matrix 3 adding FA to column 82 
	-- signal N4_6_82 : std_logic;
	-- signal N4_7_83 : std_logic;
	FA1336 : full_adder port map (N0_39_82,N0_40_82,N0_41_82,N4_6_82,N4_7_83);
-- In matrix 3 adding FA to column 82 
	-- signal N4_8_82 : std_logic;
	-- signal N4_9_83 : std_logic;
	FA1337 : full_adder port map (N0_42_82,N0_43_82,N0_44_82,N4_8_82,N4_9_83);
-- In matrix 3 adding FA to column 82 
	-- signal N4_10_82 : std_logic;
	-- signal N4_11_83 : std_logic;
	FA1338 : full_adder port map (N0_45_82,N0_46_82,N0_47_82,N4_10_82,N4_11_83);
-- In matrix 3 adding FA to column 82 
	-- signal N4_12_82 : std_logic;
	-- signal N4_13_83 : std_logic;
	FA1339 : full_adder port map (N0_48_82,N0_49_82,N0_50_82,N4_12_82,N4_13_83);
-- In matrix 3 adding FA to column 82 
	-- signal N4_14_82 : std_logic;
	-- signal N4_15_83 : std_logic;
	FA1340 : full_adder port map (N0_51_82,N0_52_82,N3_1_82,N4_14_82,N4_15_83);
-- In matrix 3 adding FA to column 83 
	-- signal N4_0_83 : std_logic;
	-- signal N4_1_84 : std_logic;
	FA1341 : full_adder port map (N0_31_83,N0_32_83,N0_33_83,N4_0_83,N4_1_84);
-- In matrix 3 adding FA to column 83 
	-- signal N4_2_83 : std_logic;
	-- signal N4_3_84 : std_logic;
	FA1342 : full_adder port map (N0_34_83,N0_35_83,N0_36_83,N4_2_83,N4_3_84);
-- In matrix 3 adding FA to column 83 
	-- signal N4_4_83 : std_logic;
	-- signal N4_5_84 : std_logic;
	FA1343 : full_adder port map (N0_37_83,N0_38_83,N0_39_83,N4_4_83,N4_5_84);
-- In matrix 3 adding FA to column 83 
	-- signal N4_6_83 : std_logic;
	-- signal N4_7_84 : std_logic;
	FA1344 : full_adder port map (N0_40_83,N0_41_83,N0_42_83,N4_6_83,N4_7_84);
-- In matrix 3 adding FA to column 83 
	-- signal N4_8_83 : std_logic;
	-- signal N4_9_84 : std_logic;
	FA1345 : full_adder port map (N0_43_83,N0_44_83,N0_45_83,N4_8_83,N4_9_84);
-- In matrix 3 adding FA to column 83 
	-- signal N4_10_83 : std_logic;
	-- signal N4_11_84 : std_logic;
	FA1346 : full_adder port map (N0_46_83,N0_47_83,N0_48_83,N4_10_83,N4_11_84);
-- In matrix 3 adding FA to column 83 
	-- signal N4_12_83 : std_logic;
	-- signal N4_13_84 : std_logic;
	FA1347 : full_adder port map (N0_49_83,N0_50_83,N0_51_83,N4_12_83,N4_13_84);
-- In matrix 3 adding FA to column 84 
	-- signal N4_0_84 : std_logic;
	-- signal N4_1_85 : std_logic;
	FA1348 : full_adder port map (N0_32_84,N0_33_84,N0_34_84,N4_0_84,N4_1_85);
-- In matrix 3 adding FA to column 84 
	-- signal N4_2_84 : std_logic;
	-- signal N4_3_85 : std_logic;
	FA1349 : full_adder port map (N0_35_84,N0_36_84,N0_37_84,N4_2_84,N4_3_85);
-- In matrix 3 adding FA to column 84 
	-- signal N4_4_84 : std_logic;
	-- signal N4_5_85 : std_logic;
	FA1350 : full_adder port map (N0_38_84,N0_39_84,N0_40_84,N4_4_84,N4_5_85);
-- In matrix 3 adding FA to column 84 
	-- signal N4_6_84 : std_logic;
	-- signal N4_7_85 : std_logic;
	FA1351 : full_adder port map (N0_41_84,N0_42_84,N0_43_84,N4_6_84,N4_7_85);
-- In matrix 3 adding FA to column 84 
	-- signal N4_8_84 : std_logic;
	-- signal N4_9_85 : std_logic;
	FA1352 : full_adder port map (N0_44_84,N0_45_84,N0_46_84,N4_8_84,N4_9_85);
-- In matrix 3 adding FA to column 84 
	-- signal N4_10_84 : std_logic;
	-- signal N4_11_85 : std_logic;
	FA1353 : full_adder port map (N0_47_84,N0_48_84,N0_49_84,N4_10_84,N4_11_85);
-- In matrix 3 adding FA to column 85 
	-- signal N4_0_85 : std_logic;
	-- signal N4_1_86 : std_logic;
	FA1354 : full_adder port map (N0_33_85,N0_34_85,N0_35_85,N4_0_85,N4_1_86);
-- In matrix 3 adding FA to column 85 
	-- signal N4_2_85 : std_logic;
	-- signal N4_3_86 : std_logic;
	FA1355 : full_adder port map (N0_36_85,N0_37_85,N0_38_85,N4_2_85,N4_3_86);
-- In matrix 3 adding FA to column 85 
	-- signal N4_4_85 : std_logic;
	-- signal N4_5_86 : std_logic;
	FA1356 : full_adder port map (N0_39_85,N0_40_85,N0_41_85,N4_4_85,N4_5_86);
-- In matrix 3 adding FA to column 85 
	-- signal N4_6_85 : std_logic;
	-- signal N4_7_86 : std_logic;
	FA1357 : full_adder port map (N0_42_85,N0_43_85,N0_44_85,N4_6_85,N4_7_86);
-- In matrix 3 adding FA to column 85 
	-- signal N4_8_85 : std_logic;
	-- signal N4_9_86 : std_logic;
	FA1358 : full_adder port map (N0_45_85,N0_46_85,N0_47_85,N4_8_85,N4_9_86);
-- In matrix 3 adding FA to column 86 
	-- signal N4_0_86 : std_logic;
	-- signal N4_1_87 : std_logic;
	FA1359 : full_adder port map (N0_34_86,N0_35_86,N0_36_86,N4_0_86,N4_1_87);
-- In matrix 3 adding FA to column 86 
	-- signal N4_2_86 : std_logic;
	-- signal N4_3_87 : std_logic;
	FA1360 : full_adder port map (N0_37_86,N0_38_86,N0_39_86,N4_2_86,N4_3_87);
-- In matrix 3 adding FA to column 86 
	-- signal N4_4_86 : std_logic;
	-- signal N4_5_87 : std_logic;
	FA1361 : full_adder port map (N0_40_86,N0_41_86,N0_42_86,N4_4_86,N4_5_87);
-- In matrix 3 adding FA to column 86 
	-- signal N4_6_86 : std_logic;
	-- signal N4_7_87 : std_logic;
	FA1362 : full_adder port map (N0_43_86,N0_44_86,N0_45_86,N4_6_86,N4_7_87);
-- In matrix 3 adding FA to column 87 
	-- signal N4_0_87 : std_logic;
	-- signal N4_1_88 : std_logic;
	FA1363 : full_adder port map (N0_35_87,N0_36_87,N0_37_87,N4_0_87,N4_1_88);
-- In matrix 3 adding FA to column 87 
	-- signal N4_2_87 : std_logic;
	-- signal N4_3_88 : std_logic;
	FA1364 : full_adder port map (N0_38_87,N0_39_87,N0_40_87,N4_2_87,N4_3_88);
-- In matrix 3 adding FA to column 87 
	-- signal N4_4_87 : std_logic;
	-- signal N4_5_88 : std_logic;
	FA1365 : full_adder port map (N0_41_87,N0_42_87,N0_43_87,N4_4_87,N4_5_88);
-- In matrix 3 adding FA to column 88 
	-- signal N4_0_88 : std_logic;
	-- signal N4_1_89 : std_logic;
	FA1366 : full_adder port map (N0_36_88,N0_37_88,N0_38_88,N4_0_88,N4_1_89);
-- In matrix 3 adding FA to column 88 
	-- signal N4_2_88 : std_logic;
	-- signal N4_3_89 : std_logic;
	FA1367 : full_adder port map (N0_39_88,N0_40_88,N0_41_88,N4_2_88,N4_3_89);
-- In matrix 3 adding FA to column 89 
	-- signal N4_0_89 : std_logic;
	-- signal N4_1_90 : std_logic;
	FA1368 : full_adder port map (N0_37_89,N0_38_89,N0_39_89,N4_0_89,N4_1_90);
	-- Elements from matrix 4 
-- In matrix 4 adding HA to column 11 
	-- signal N5_0_11 : std_logic;
	-- signal N5_1_12 : std_logic;
	HA39 : half_adder port map (N0_0_11,N0_1_11,N5_0_11,N5_1_12);
-- In matrix 4 adding FA to column 12 
	-- signal N5_0_12 : std_logic;
	-- signal N5_1_13 : std_logic;
	FA1369 : full_adder port map (N0_0_12,N0_1_12,N0_2_12,N5_0_12,N5_1_13);
-- In matrix 4 adding HA to column 12 
	-- signal N5_2_12 : std_logic;
	-- signal N5_3_13 : std_logic;
	HA40 : half_adder port map (N0_3_12,N0_4_12,N5_2_12,N5_3_13);
-- In matrix 4 adding FA to column 13 
	-- signal N5_0_13 : std_logic;
	-- signal N5_1_14 : std_logic;
	FA1370 : full_adder port map (N0_0_13,N0_1_13,N0_2_13,N5_0_13,N5_1_14);
-- In matrix 4 adding FA to column 13 
	-- signal N5_2_13 : std_logic;
	-- signal N5_3_14 : std_logic;
	FA1371 : full_adder port map (N0_3_13,N0_4_13,N0_5_13,N5_2_13,N5_3_14);
-- In matrix 4 adding HA to column 13 
	-- signal N5_4_13 : std_logic;
	-- signal N5_5_14 : std_logic;
	HA41 : half_adder port map (N0_6_13,N0_7_13,N5_4_13,N5_5_14);
-- In matrix 4 adding FA to column 14 
	-- signal N5_0_14 : std_logic;
	-- signal N5_1_15 : std_logic;
	FA1372 : full_adder port map (N0_0_14,N0_1_14,N0_2_14,N5_0_14,N5_1_15);
-- In matrix 4 adding FA to column 14 
	-- signal N5_2_14 : std_logic;
	-- signal N5_3_15 : std_logic;
	FA1373 : full_adder port map (N0_3_14,N0_4_14,N0_5_14,N5_2_14,N5_3_15);
-- In matrix 4 adding FA to column 14 
	-- signal N5_4_14 : std_logic;
	-- signal N5_5_15 : std_logic;
	FA1374 : full_adder port map (N0_6_14,N0_7_14,N0_8_14,N5_4_14,N5_5_15);
-- In matrix 4 adding HA to column 14 
	-- signal N5_6_14 : std_logic;
	-- signal N5_7_15 : std_logic;
	HA42 : half_adder port map (N0_9_14,N0_10_14,N5_6_14,N5_7_15);
-- In matrix 4 adding FA to column 15 
	-- signal N5_0_15 : std_logic;
	-- signal N5_1_16 : std_logic;
	FA1375 : full_adder port map (N0_0_15,N0_1_15,N0_2_15,N5_0_15,N5_1_16);
-- In matrix 4 adding FA to column 15 
	-- signal N5_2_15 : std_logic;
	-- signal N5_3_16 : std_logic;
	FA1376 : full_adder port map (N0_3_15,N0_4_15,N0_5_15,N5_2_15,N5_3_16);
-- In matrix 4 adding FA to column 15 
	-- signal N5_4_15 : std_logic;
	-- signal N5_5_16 : std_logic;
	FA1377 : full_adder port map (N0_6_15,N0_7_15,N0_8_15,N5_4_15,N5_5_16);
-- In matrix 4 adding FA to column 15 
	-- signal N5_6_15 : std_logic;
	-- signal N5_7_16 : std_logic;
	FA1378 : full_adder port map (N0_9_15,N0_10_15,N0_11_15,N5_6_15,N5_7_16);
-- In matrix 4 adding HA to column 15 
	-- signal N5_8_15 : std_logic;
	-- signal N5_9_16 : std_logic;
	HA43 : half_adder port map (N0_12_15,N0_13_15,N5_8_15,N5_9_16);
-- In matrix 4 adding FA to column 16 
	-- signal N5_0_16 : std_logic;
	-- signal N5_1_17 : std_logic;
	FA1379 : full_adder port map (N0_2_16,N0_3_16,N0_4_16,N5_0_16,N5_1_17);
-- In matrix 4 adding FA to column 16 
	-- signal N5_2_16 : std_logic;
	-- signal N5_3_17 : std_logic;
	FA1380 : full_adder port map (N0_5_16,N0_6_16,N0_7_16,N5_2_16,N5_3_17);
-- In matrix 4 adding FA to column 16 
	-- signal N5_4_16 : std_logic;
	-- signal N5_5_17 : std_logic;
	FA1381 : full_adder port map (N0_8_16,N0_9_16,N0_10_16,N5_4_16,N5_5_17);
-- In matrix 4 adding FA to column 16 
	-- signal N5_6_16 : std_logic;
	-- signal N5_7_17 : std_logic;
	FA1382 : full_adder port map (N0_11_16,N0_12_16,N0_13_16,N5_6_16,N5_7_17);
-- In matrix 4 adding FA to column 16 
	-- signal N5_8_16 : std_logic;
	-- signal N5_9_17 : std_logic;
	FA1383 : full_adder port map (N0_14_16,N0_15_16,N0_16_16,N5_8_16,N5_9_17);
-- In matrix 4 adding FA to column 17 
	-- signal N5_0_17 : std_logic;
	-- signal N5_1_18 : std_logic;
	FA1384 : full_adder port map (N0_5_17,N0_6_17,N0_7_17,N5_0_17,N5_1_18);
-- In matrix 4 adding FA to column 17 
	-- signal N5_2_17 : std_logic;
	-- signal N5_3_18 : std_logic;
	FA1385 : full_adder port map (N0_8_17,N0_9_17,N0_10_17,N5_2_17,N5_3_18);
-- In matrix 4 adding FA to column 17 
	-- signal N5_4_17 : std_logic;
	-- signal N5_5_18 : std_logic;
	FA1386 : full_adder port map (N0_11_17,N0_12_17,N0_13_17,N5_4_17,N5_5_18);
-- In matrix 4 adding FA to column 17 
	-- signal N5_6_17 : std_logic;
	-- signal N5_7_18 : std_logic;
	FA1387 : full_adder port map (N0_14_17,N0_15_17,N0_16_17,N5_6_17,N5_7_18);
-- In matrix 4 adding FA to column 17 
	-- signal N5_8_17 : std_logic;
	-- signal N5_9_18 : std_logic;
	FA1388 : full_adder port map (N0_17_17,N4_0_17,N4_1_17,N5_8_17,N5_9_18);
-- In matrix 4 adding FA to column 18 
	-- signal N5_0_18 : std_logic;
	-- signal N5_1_19 : std_logic;
	FA1389 : full_adder port map (N0_8_18,N0_9_18,N0_10_18,N5_0_18,N5_1_19);
-- In matrix 4 adding FA to column 18 
	-- signal N5_2_18 : std_logic;
	-- signal N5_3_19 : std_logic;
	FA1390 : full_adder port map (N0_11_18,N0_12_18,N0_13_18,N5_2_18,N5_3_19);
-- In matrix 4 adding FA to column 18 
	-- signal N5_4_18 : std_logic;
	-- signal N5_5_19 : std_logic;
	FA1391 : full_adder port map (N0_14_18,N0_15_18,N0_16_18,N5_4_18,N5_5_19);
-- In matrix 4 adding FA to column 18 
	-- signal N5_6_18 : std_logic;
	-- signal N5_7_19 : std_logic;
	FA1392 : full_adder port map (N0_17_18,N0_18_18,N4_0_18,N5_6_18,N5_7_19);
-- In matrix 4 adding FA to column 18 
	-- signal N5_8_18 : std_logic;
	-- signal N5_9_19 : std_logic;
	FA1393 : full_adder port map (N4_1_18,N4_2_18,N4_3_18,N5_8_18,N5_9_19);
-- In matrix 4 adding FA to column 19 
	-- signal N5_0_19 : std_logic;
	-- signal N5_1_20 : std_logic;
	FA1394 : full_adder port map (N0_11_19,N0_12_19,N0_13_19,N5_0_19,N5_1_20);
-- In matrix 4 adding FA to column 19 
	-- signal N5_2_19 : std_logic;
	-- signal N5_3_20 : std_logic;
	FA1395 : full_adder port map (N0_14_19,N0_15_19,N0_16_19,N5_2_19,N5_3_20);
-- In matrix 4 adding FA to column 19 
	-- signal N5_4_19 : std_logic;
	-- signal N5_5_20 : std_logic;
	FA1396 : full_adder port map (N0_17_19,N0_18_19,N0_19_19,N5_4_19,N5_5_20);
-- In matrix 4 adding FA to column 19 
	-- signal N5_6_19 : std_logic;
	-- signal N5_7_20 : std_logic;
	FA1397 : full_adder port map (N4_0_19,N4_1_19,N4_2_19,N5_6_19,N5_7_20);
-- In matrix 4 adding FA to column 19 
	-- signal N5_8_19 : std_logic;
	-- signal N5_9_20 : std_logic;
	FA1398 : full_adder port map (N4_3_19,N4_4_19,N4_5_19,N5_8_19,N5_9_20);
-- In matrix 4 adding FA to column 20 
	-- signal N5_0_20 : std_logic;
	-- signal N5_1_21 : std_logic;
	FA1399 : full_adder port map (N0_14_20,N0_15_20,N0_16_20,N5_0_20,N5_1_21);
-- In matrix 4 adding FA to column 20 
	-- signal N5_2_20 : std_logic;
	-- signal N5_3_21 : std_logic;
	FA1400 : full_adder port map (N0_17_20,N0_18_20,N0_19_20,N5_2_20,N5_3_21);
-- In matrix 4 adding FA to column 20 
	-- signal N5_4_20 : std_logic;
	-- signal N5_5_21 : std_logic;
	FA1401 : full_adder port map (N0_20_20,N4_0_20,N4_1_20,N5_4_20,N5_5_21);
-- In matrix 4 adding FA to column 20 
	-- signal N5_6_20 : std_logic;
	-- signal N5_7_21 : std_logic;
	FA1402 : full_adder port map (N4_2_20,N4_3_20,N4_4_20,N5_6_20,N5_7_21);
-- In matrix 4 adding FA to column 20 
	-- signal N5_8_20 : std_logic;
	-- signal N5_9_21 : std_logic;
	FA1403 : full_adder port map (N4_5_20,N4_6_20,N4_7_20,N5_8_20,N5_9_21);
-- In matrix 4 adding FA to column 21 
	-- signal N5_0_21 : std_logic;
	-- signal N5_1_22 : std_logic;
	FA1404 : full_adder port map (N0_17_21,N0_18_21,N0_19_21,N5_0_21,N5_1_22);
-- In matrix 4 adding FA to column 21 
	-- signal N5_2_21 : std_logic;
	-- signal N5_3_22 : std_logic;
	FA1405 : full_adder port map (N0_20_21,N0_21_21,N4_0_21,N5_2_21,N5_3_22);
-- In matrix 4 adding FA to column 21 
	-- signal N5_4_21 : std_logic;
	-- signal N5_5_22 : std_logic;
	FA1406 : full_adder port map (N4_1_21,N4_2_21,N4_3_21,N5_4_21,N5_5_22);
-- In matrix 4 adding FA to column 21 
	-- signal N5_6_21 : std_logic;
	-- signal N5_7_22 : std_logic;
	FA1407 : full_adder port map (N4_4_21,N4_5_21,N4_6_21,N5_6_21,N5_7_22);
-- In matrix 4 adding FA to column 21 
	-- signal N5_8_21 : std_logic;
	-- signal N5_9_22 : std_logic;
	FA1408 : full_adder port map (N4_7_21,N4_8_21,N4_9_21,N5_8_21,N5_9_22);
-- In matrix 4 adding FA to column 22 
	-- signal N5_0_22 : std_logic;
	-- signal N5_1_23 : std_logic;
	FA1409 : full_adder port map (N0_20_22,N0_21_22,N0_22_22,N5_0_22,N5_1_23);
-- In matrix 4 adding FA to column 22 
	-- signal N5_2_22 : std_logic;
	-- signal N5_3_23 : std_logic;
	FA1410 : full_adder port map (N4_0_22,N4_1_22,N4_2_22,N5_2_22,N5_3_23);
-- In matrix 4 adding FA to column 22 
	-- signal N5_4_22 : std_logic;
	-- signal N5_5_23 : std_logic;
	FA1411 : full_adder port map (N4_3_22,N4_4_22,N4_5_22,N5_4_22,N5_5_23);
-- In matrix 4 adding FA to column 22 
	-- signal N5_6_22 : std_logic;
	-- signal N5_7_23 : std_logic;
	FA1412 : full_adder port map (N4_6_22,N4_7_22,N4_8_22,N5_6_22,N5_7_23);
-- In matrix 4 adding FA to column 22 
	-- signal N5_8_22 : std_logic;
	-- signal N5_9_23 : std_logic;
	FA1413 : full_adder port map (N4_9_22,N4_10_22,N4_11_22,N5_8_22,N5_9_23);
-- In matrix 4 adding FA to column 23 
	-- signal N5_0_23 : std_logic;
	-- signal N5_1_24 : std_logic;
	FA1414 : full_adder port map (N0_23_23,N4_0_23,N4_1_23,N5_0_23,N5_1_24);
-- In matrix 4 adding FA to column 23 
	-- signal N5_2_23 : std_logic;
	-- signal N5_3_24 : std_logic;
	FA1415 : full_adder port map (N4_2_23,N4_3_23,N4_4_23,N5_2_23,N5_3_24);
-- In matrix 4 adding FA to column 23 
	-- signal N5_4_23 : std_logic;
	-- signal N5_5_24 : std_logic;
	FA1416 : full_adder port map (N4_5_23,N4_6_23,N4_7_23,N5_4_23,N5_5_24);
-- In matrix 4 adding FA to column 23 
	-- signal N5_6_23 : std_logic;
	-- signal N5_7_24 : std_logic;
	FA1417 : full_adder port map (N4_8_23,N4_9_23,N4_10_23,N5_6_23,N5_7_24);
-- In matrix 4 adding FA to column 23 
	-- signal N5_8_23 : std_logic;
	-- signal N5_9_24 : std_logic;
	FA1418 : full_adder port map (N4_11_23,N4_12_23,N4_13_23,N5_8_23,N5_9_24);
-- In matrix 4 adding FA to column 24 
	-- signal N5_0_24 : std_logic;
	-- signal N5_1_25 : std_logic;
	FA1419 : full_adder port map (N4_0_24,N4_1_24,N4_2_24,N5_0_24,N5_1_25);
-- In matrix 4 adding FA to column 24 
	-- signal N5_2_24 : std_logic;
	-- signal N5_3_25 : std_logic;
	FA1420 : full_adder port map (N4_3_24,N4_4_24,N4_5_24,N5_2_24,N5_3_25);
-- In matrix 4 adding FA to column 24 
	-- signal N5_4_24 : std_logic;
	-- signal N5_5_25 : std_logic;
	FA1421 : full_adder port map (N4_6_24,N4_7_24,N4_8_24,N5_4_24,N5_5_25);
-- In matrix 4 adding FA to column 24 
	-- signal N5_6_24 : std_logic;
	-- signal N5_7_25 : std_logic;
	FA1422 : full_adder port map (N4_9_24,N4_10_24,N4_11_24,N5_6_24,N5_7_25);
-- In matrix 4 adding FA to column 24 
	-- signal N5_8_24 : std_logic;
	-- signal N5_9_25 : std_logic;
	FA1423 : full_adder port map (N4_12_24,N4_13_24,N4_14_24,N5_8_24,N5_9_25);
-- In matrix 4 adding FA to column 25 
	-- signal N5_0_25 : std_logic;
	-- signal N5_1_26 : std_logic;
	FA1424 : full_adder port map (N4_0_25,N4_1_25,N4_2_25,N5_0_25,N5_1_26);
-- In matrix 4 adding FA to column 25 
	-- signal N5_2_25 : std_logic;
	-- signal N5_3_26 : std_logic;
	FA1425 : full_adder port map (N4_3_25,N4_4_25,N4_5_25,N5_2_25,N5_3_26);
-- In matrix 4 adding FA to column 25 
	-- signal N5_4_25 : std_logic;
	-- signal N5_5_26 : std_logic;
	FA1426 : full_adder port map (N4_6_25,N4_7_25,N4_8_25,N5_4_25,N5_5_26);
-- In matrix 4 adding FA to column 25 
	-- signal N5_6_25 : std_logic;
	-- signal N5_7_26 : std_logic;
	FA1427 : full_adder port map (N4_9_25,N4_10_25,N4_11_25,N5_6_25,N5_7_26);
-- In matrix 4 adding FA to column 25 
	-- signal N5_8_25 : std_logic;
	-- signal N5_9_26 : std_logic;
	FA1428 : full_adder port map (N4_12_25,N4_13_25,N4_14_25,N5_8_25,N5_9_26);
-- In matrix 4 adding FA to column 26 
	-- signal N5_0_26 : std_logic;
	-- signal N5_1_27 : std_logic;
	FA1429 : full_adder port map (N4_0_26,N4_1_26,N4_2_26,N5_0_26,N5_1_27);
-- In matrix 4 adding FA to column 26 
	-- signal N5_2_26 : std_logic;
	-- signal N5_3_27 : std_logic;
	FA1430 : full_adder port map (N4_3_26,N4_4_26,N4_5_26,N5_2_26,N5_3_27);
-- In matrix 4 adding FA to column 26 
	-- signal N5_4_26 : std_logic;
	-- signal N5_5_27 : std_logic;
	FA1431 : full_adder port map (N4_6_26,N4_7_26,N4_8_26,N5_4_26,N5_5_27);
-- In matrix 4 adding FA to column 26 
	-- signal N5_6_26 : std_logic;
	-- signal N5_7_27 : std_logic;
	FA1432 : full_adder port map (N4_9_26,N4_10_26,N4_11_26,N5_6_26,N5_7_27);
-- In matrix 4 adding FA to column 26 
	-- signal N5_8_26 : std_logic;
	-- signal N5_9_27 : std_logic;
	FA1433 : full_adder port map (N4_12_26,N4_13_26,N4_14_26,N5_8_26,N5_9_27);
-- In matrix 4 adding FA to column 27 
	-- signal N5_0_27 : std_logic;
	-- signal N5_1_28 : std_logic;
	FA1434 : full_adder port map (N4_0_27,N4_1_27,N4_2_27,N5_0_27,N5_1_28);
-- In matrix 4 adding FA to column 27 
	-- signal N5_2_27 : std_logic;
	-- signal N5_3_28 : std_logic;
	FA1435 : full_adder port map (N4_3_27,N4_4_27,N4_5_27,N5_2_27,N5_3_28);
-- In matrix 4 adding FA to column 27 
	-- signal N5_4_27 : std_logic;
	-- signal N5_5_28 : std_logic;
	FA1436 : full_adder port map (N4_6_27,N4_7_27,N4_8_27,N5_4_27,N5_5_28);
-- In matrix 4 adding FA to column 27 
	-- signal N5_6_27 : std_logic;
	-- signal N5_7_28 : std_logic;
	FA1437 : full_adder port map (N4_9_27,N4_10_27,N4_11_27,N5_6_27,N5_7_28);
-- In matrix 4 adding FA to column 27 
	-- signal N5_8_27 : std_logic;
	-- signal N5_9_28 : std_logic;
	FA1438 : full_adder port map (N4_12_27,N4_13_27,N4_14_27,N5_8_27,N5_9_28);
-- In matrix 4 adding FA to column 28 
	-- signal N5_0_28 : std_logic;
	-- signal N5_1_29 : std_logic;
	FA1439 : full_adder port map (N4_0_28,N4_1_28,N4_2_28,N5_0_28,N5_1_29);
-- In matrix 4 adding FA to column 28 
	-- signal N5_2_28 : std_logic;
	-- signal N5_3_29 : std_logic;
	FA1440 : full_adder port map (N4_3_28,N4_4_28,N4_5_28,N5_2_28,N5_3_29);
-- In matrix 4 adding FA to column 28 
	-- signal N5_4_28 : std_logic;
	-- signal N5_5_29 : std_logic;
	FA1441 : full_adder port map (N4_6_28,N4_7_28,N4_8_28,N5_4_28,N5_5_29);
-- In matrix 4 adding FA to column 28 
	-- signal N5_6_28 : std_logic;
	-- signal N5_7_29 : std_logic;
	FA1442 : full_adder port map (N4_9_28,N4_10_28,N4_11_28,N5_6_28,N5_7_29);
-- In matrix 4 adding FA to column 28 
	-- signal N5_8_28 : std_logic;
	-- signal N5_9_29 : std_logic;
	FA1443 : full_adder port map (N4_12_28,N4_13_28,N4_14_28,N5_8_28,N5_9_29);
-- In matrix 4 adding FA to column 29 
	-- signal N5_0_29 : std_logic;
	-- signal N5_1_30 : std_logic;
	FA1444 : full_adder port map (N4_0_29,N4_1_29,N4_2_29,N5_0_29,N5_1_30);
-- In matrix 4 adding FA to column 29 
	-- signal N5_2_29 : std_logic;
	-- signal N5_3_30 : std_logic;
	FA1445 : full_adder port map (N4_3_29,N4_4_29,N4_5_29,N5_2_29,N5_3_30);
-- In matrix 4 adding FA to column 29 
	-- signal N5_4_29 : std_logic;
	-- signal N5_5_30 : std_logic;
	FA1446 : full_adder port map (N4_6_29,N4_7_29,N4_8_29,N5_4_29,N5_5_30);
-- In matrix 4 adding FA to column 29 
	-- signal N5_6_29 : std_logic;
	-- signal N5_7_30 : std_logic;
	FA1447 : full_adder port map (N4_9_29,N4_10_29,N4_11_29,N5_6_29,N5_7_30);
-- In matrix 4 adding FA to column 29 
	-- signal N5_8_29 : std_logic;
	-- signal N5_9_30 : std_logic;
	FA1448 : full_adder port map (N4_12_29,N4_13_29,N4_14_29,N5_8_29,N5_9_30);
-- In matrix 4 adding FA to column 30 
	-- signal N5_0_30 : std_logic;
	-- signal N5_1_31 : std_logic;
	FA1449 : full_adder port map (N4_0_30,N4_1_30,N4_2_30,N5_0_30,N5_1_31);
-- In matrix 4 adding FA to column 30 
	-- signal N5_2_30 : std_logic;
	-- signal N5_3_31 : std_logic;
	FA1450 : full_adder port map (N4_3_30,N4_4_30,N4_5_30,N5_2_30,N5_3_31);
-- In matrix 4 adding FA to column 30 
	-- signal N5_4_30 : std_logic;
	-- signal N5_5_31 : std_logic;
	FA1451 : full_adder port map (N4_6_30,N4_7_30,N4_8_30,N5_4_30,N5_5_31);
-- In matrix 4 adding FA to column 30 
	-- signal N5_6_30 : std_logic;
	-- signal N5_7_31 : std_logic;
	FA1452 : full_adder port map (N4_9_30,N4_10_30,N4_11_30,N5_6_30,N5_7_31);
-- In matrix 4 adding FA to column 30 
	-- signal N5_8_30 : std_logic;
	-- signal N5_9_31 : std_logic;
	FA1453 : full_adder port map (N4_12_30,N4_13_30,N4_14_30,N5_8_30,N5_9_31);
-- In matrix 4 adding FA to column 31 
	-- signal N5_0_31 : std_logic;
	-- signal N5_1_32 : std_logic;
	FA1454 : full_adder port map (N4_0_31,N4_1_31,N4_2_31,N5_0_31,N5_1_32);
-- In matrix 4 adding FA to column 31 
	-- signal N5_2_31 : std_logic;
	-- signal N5_3_32 : std_logic;
	FA1455 : full_adder port map (N4_3_31,N4_4_31,N4_5_31,N5_2_31,N5_3_32);
-- In matrix 4 adding FA to column 31 
	-- signal N5_4_31 : std_logic;
	-- signal N5_5_32 : std_logic;
	FA1456 : full_adder port map (N4_6_31,N4_7_31,N4_8_31,N5_4_31,N5_5_32);
-- In matrix 4 adding FA to column 31 
	-- signal N5_6_31 : std_logic;
	-- signal N5_7_32 : std_logic;
	FA1457 : full_adder port map (N4_9_31,N4_10_31,N4_11_31,N5_6_31,N5_7_32);
-- In matrix 4 adding FA to column 31 
	-- signal N5_8_31 : std_logic;
	-- signal N5_9_32 : std_logic;
	FA1458 : full_adder port map (N4_12_31,N4_13_31,N4_14_31,N5_8_31,N5_9_32);
-- In matrix 4 adding FA to column 32 
	-- signal N5_0_32 : std_logic;
	-- signal N5_1_33 : std_logic;
	FA1459 : full_adder port map (N4_0_32,N4_1_32,N4_2_32,N5_0_32,N5_1_33);
-- In matrix 4 adding FA to column 32 
	-- signal N5_2_32 : std_logic;
	-- signal N5_3_33 : std_logic;
	FA1460 : full_adder port map (N4_3_32,N4_4_32,N4_5_32,N5_2_32,N5_3_33);
-- In matrix 4 adding FA to column 32 
	-- signal N5_4_32 : std_logic;
	-- signal N5_5_33 : std_logic;
	FA1461 : full_adder port map (N4_6_32,N4_7_32,N4_8_32,N5_4_32,N5_5_33);
-- In matrix 4 adding FA to column 32 
	-- signal N5_6_32 : std_logic;
	-- signal N5_7_33 : std_logic;
	FA1462 : full_adder port map (N4_9_32,N4_10_32,N4_11_32,N5_6_32,N5_7_33);
-- In matrix 4 adding FA to column 32 
	-- signal N5_8_32 : std_logic;
	-- signal N5_9_33 : std_logic;
	FA1463 : full_adder port map (N4_12_32,N4_13_32,N4_14_32,N5_8_32,N5_9_33);
-- In matrix 4 adding FA to column 33 
	-- signal N5_0_33 : std_logic;
	-- signal N5_1_34 : std_logic;
	FA1464 : full_adder port map (N4_0_33,N4_1_33,N4_2_33,N5_0_33,N5_1_34);
-- In matrix 4 adding FA to column 33 
	-- signal N5_2_33 : std_logic;
	-- signal N5_3_34 : std_logic;
	FA1465 : full_adder port map (N4_3_33,N4_4_33,N4_5_33,N5_2_33,N5_3_34);
-- In matrix 4 adding FA to column 33 
	-- signal N5_4_33 : std_logic;
	-- signal N5_5_34 : std_logic;
	FA1466 : full_adder port map (N4_6_33,N4_7_33,N4_8_33,N5_4_33,N5_5_34);
-- In matrix 4 adding FA to column 33 
	-- signal N5_6_33 : std_logic;
	-- signal N5_7_34 : std_logic;
	FA1467 : full_adder port map (N4_9_33,N4_10_33,N4_11_33,N5_6_33,N5_7_34);
-- In matrix 4 adding FA to column 33 
	-- signal N5_8_33 : std_logic;
	-- signal N5_9_34 : std_logic;
	FA1468 : full_adder port map (N4_12_33,N4_13_33,N4_14_33,N5_8_33,N5_9_34);
-- In matrix 4 adding FA to column 34 
	-- signal N5_0_34 : std_logic;
	-- signal N5_1_35 : std_logic;
	FA1469 : full_adder port map (N4_0_34,N4_1_34,N4_2_34,N5_0_34,N5_1_35);
-- In matrix 4 adding FA to column 34 
	-- signal N5_2_34 : std_logic;
	-- signal N5_3_35 : std_logic;
	FA1470 : full_adder port map (N4_3_34,N4_4_34,N4_5_34,N5_2_34,N5_3_35);
-- In matrix 4 adding FA to column 34 
	-- signal N5_4_34 : std_logic;
	-- signal N5_5_35 : std_logic;
	FA1471 : full_adder port map (N4_6_34,N4_7_34,N4_8_34,N5_4_34,N5_5_35);
-- In matrix 4 adding FA to column 34 
	-- signal N5_6_34 : std_logic;
	-- signal N5_7_35 : std_logic;
	FA1472 : full_adder port map (N4_9_34,N4_10_34,N4_11_34,N5_6_34,N5_7_35);
-- In matrix 4 adding FA to column 34 
	-- signal N5_8_34 : std_logic;
	-- signal N5_9_35 : std_logic;
	FA1473 : full_adder port map (N4_12_34,N4_13_34,N4_14_34,N5_8_34,N5_9_35);
-- In matrix 4 adding FA to column 35 
	-- signal N5_0_35 : std_logic;
	-- signal N5_1_36 : std_logic;
	FA1474 : full_adder port map (N4_0_35,N4_1_35,N4_2_35,N5_0_35,N5_1_36);
-- In matrix 4 adding FA to column 35 
	-- signal N5_2_35 : std_logic;
	-- signal N5_3_36 : std_logic;
	FA1475 : full_adder port map (N4_3_35,N4_4_35,N4_5_35,N5_2_35,N5_3_36);
-- In matrix 4 adding FA to column 35 
	-- signal N5_4_35 : std_logic;
	-- signal N5_5_36 : std_logic;
	FA1476 : full_adder port map (N4_6_35,N4_7_35,N4_8_35,N5_4_35,N5_5_36);
-- In matrix 4 adding FA to column 35 
	-- signal N5_6_35 : std_logic;
	-- signal N5_7_36 : std_logic;
	FA1477 : full_adder port map (N4_9_35,N4_10_35,N4_11_35,N5_6_35,N5_7_36);
-- In matrix 4 adding FA to column 35 
	-- signal N5_8_35 : std_logic;
	-- signal N5_9_36 : std_logic;
	FA1478 : full_adder port map (N4_12_35,N4_13_35,N4_14_35,N5_8_35,N5_9_36);
-- In matrix 4 adding FA to column 36 
	-- signal N5_0_36 : std_logic;
	-- signal N5_1_37 : std_logic;
	FA1479 : full_adder port map (N4_0_36,N4_1_36,N4_2_36,N5_0_36,N5_1_37);
-- In matrix 4 adding FA to column 36 
	-- signal N5_2_36 : std_logic;
	-- signal N5_3_37 : std_logic;
	FA1480 : full_adder port map (N4_3_36,N4_4_36,N4_5_36,N5_2_36,N5_3_37);
-- In matrix 4 adding FA to column 36 
	-- signal N5_4_36 : std_logic;
	-- signal N5_5_37 : std_logic;
	FA1481 : full_adder port map (N4_6_36,N4_7_36,N4_8_36,N5_4_36,N5_5_37);
-- In matrix 4 adding FA to column 36 
	-- signal N5_6_36 : std_logic;
	-- signal N5_7_37 : std_logic;
	FA1482 : full_adder port map (N4_9_36,N4_10_36,N4_11_36,N5_6_36,N5_7_37);
-- In matrix 4 adding FA to column 36 
	-- signal N5_8_36 : std_logic;
	-- signal N5_9_37 : std_logic;
	FA1483 : full_adder port map (N4_12_36,N4_13_36,N4_14_36,N5_8_36,N5_9_37);
-- In matrix 4 adding FA to column 37 
	-- signal N5_0_37 : std_logic;
	-- signal N5_1_38 : std_logic;
	FA1484 : full_adder port map (N4_0_37,N4_1_37,N4_2_37,N5_0_37,N5_1_38);
-- In matrix 4 adding FA to column 37 
	-- signal N5_2_37 : std_logic;
	-- signal N5_3_38 : std_logic;
	FA1485 : full_adder port map (N4_3_37,N4_4_37,N4_5_37,N5_2_37,N5_3_38);
-- In matrix 4 adding FA to column 37 
	-- signal N5_4_37 : std_logic;
	-- signal N5_5_38 : std_logic;
	FA1486 : full_adder port map (N4_6_37,N4_7_37,N4_8_37,N5_4_37,N5_5_38);
-- In matrix 4 adding FA to column 37 
	-- signal N5_6_37 : std_logic;
	-- signal N5_7_38 : std_logic;
	FA1487 : full_adder port map (N4_9_37,N4_10_37,N4_11_37,N5_6_37,N5_7_38);
-- In matrix 4 adding FA to column 37 
	-- signal N5_8_37 : std_logic;
	-- signal N5_9_38 : std_logic;
	FA1488 : full_adder port map (N4_12_37,N4_13_37,N4_14_37,N5_8_37,N5_9_38);
-- In matrix 4 adding FA to column 38 
	-- signal N5_0_38 : std_logic;
	-- signal N5_1_39 : std_logic;
	FA1489 : full_adder port map (N4_0_38,N4_1_38,N4_2_38,N5_0_38,N5_1_39);
-- In matrix 4 adding FA to column 38 
	-- signal N5_2_38 : std_logic;
	-- signal N5_3_39 : std_logic;
	FA1490 : full_adder port map (N4_3_38,N4_4_38,N4_5_38,N5_2_38,N5_3_39);
-- In matrix 4 adding FA to column 38 
	-- signal N5_4_38 : std_logic;
	-- signal N5_5_39 : std_logic;
	FA1491 : full_adder port map (N4_6_38,N4_7_38,N4_8_38,N5_4_38,N5_5_39);
-- In matrix 4 adding FA to column 38 
	-- signal N5_6_38 : std_logic;
	-- signal N5_7_39 : std_logic;
	FA1492 : full_adder port map (N4_9_38,N4_10_38,N4_11_38,N5_6_38,N5_7_39);
-- In matrix 4 adding FA to column 38 
	-- signal N5_8_38 : std_logic;
	-- signal N5_9_39 : std_logic;
	FA1493 : full_adder port map (N4_12_38,N4_13_38,N4_14_38,N5_8_38,N5_9_39);
-- In matrix 4 adding FA to column 39 
	-- signal N5_0_39 : std_logic;
	-- signal N5_1_40 : std_logic;
	FA1494 : full_adder port map (N4_0_39,N4_1_39,N4_2_39,N5_0_39,N5_1_40);
-- In matrix 4 adding FA to column 39 
	-- signal N5_2_39 : std_logic;
	-- signal N5_3_40 : std_logic;
	FA1495 : full_adder port map (N4_3_39,N4_4_39,N4_5_39,N5_2_39,N5_3_40);
-- In matrix 4 adding FA to column 39 
	-- signal N5_4_39 : std_logic;
	-- signal N5_5_40 : std_logic;
	FA1496 : full_adder port map (N4_6_39,N4_7_39,N4_8_39,N5_4_39,N5_5_40);
-- In matrix 4 adding FA to column 39 
	-- signal N5_6_39 : std_logic;
	-- signal N5_7_40 : std_logic;
	FA1497 : full_adder port map (N4_9_39,N4_10_39,N4_11_39,N5_6_39,N5_7_40);
-- In matrix 4 adding FA to column 39 
	-- signal N5_8_39 : std_logic;
	-- signal N5_9_40 : std_logic;
	FA1498 : full_adder port map (N4_12_39,N4_13_39,N4_14_39,N5_8_39,N5_9_40);
-- In matrix 4 adding FA to column 40 
	-- signal N5_0_40 : std_logic;
	-- signal N5_1_41 : std_logic;
	FA1499 : full_adder port map (N4_0_40,N4_1_40,N4_2_40,N5_0_40,N5_1_41);
-- In matrix 4 adding FA to column 40 
	-- signal N5_2_40 : std_logic;
	-- signal N5_3_41 : std_logic;
	FA1500 : full_adder port map (N4_3_40,N4_4_40,N4_5_40,N5_2_40,N5_3_41);
-- In matrix 4 adding FA to column 40 
	-- signal N5_4_40 : std_logic;
	-- signal N5_5_41 : std_logic;
	FA1501 : full_adder port map (N4_6_40,N4_7_40,N4_8_40,N5_4_40,N5_5_41);
-- In matrix 4 adding FA to column 40 
	-- signal N5_6_40 : std_logic;
	-- signal N5_7_41 : std_logic;
	FA1502 : full_adder port map (N4_9_40,N4_10_40,N4_11_40,N5_6_40,N5_7_41);
-- In matrix 4 adding FA to column 40 
	-- signal N5_8_40 : std_logic;
	-- signal N5_9_41 : std_logic;
	FA1503 : full_adder port map (N4_12_40,N4_13_40,N4_14_40,N5_8_40,N5_9_41);
-- In matrix 4 adding FA to column 41 
	-- signal N5_0_41 : std_logic;
	-- signal N5_1_42 : std_logic;
	FA1504 : full_adder port map (N4_0_41,N4_1_41,N4_2_41,N5_0_41,N5_1_42);
-- In matrix 4 adding FA to column 41 
	-- signal N5_2_41 : std_logic;
	-- signal N5_3_42 : std_logic;
	FA1505 : full_adder port map (N4_3_41,N4_4_41,N4_5_41,N5_2_41,N5_3_42);
-- In matrix 4 adding FA to column 41 
	-- signal N5_4_41 : std_logic;
	-- signal N5_5_42 : std_logic;
	FA1506 : full_adder port map (N4_6_41,N4_7_41,N4_8_41,N5_4_41,N5_5_42);
-- In matrix 4 adding FA to column 41 
	-- signal N5_6_41 : std_logic;
	-- signal N5_7_42 : std_logic;
	FA1507 : full_adder port map (N4_9_41,N4_10_41,N4_11_41,N5_6_41,N5_7_42);
-- In matrix 4 adding FA to column 41 
	-- signal N5_8_41 : std_logic;
	-- signal N5_9_42 : std_logic;
	FA1508 : full_adder port map (N4_12_41,N4_13_41,N4_14_41,N5_8_41,N5_9_42);
-- In matrix 4 adding FA to column 42 
	-- signal N5_0_42 : std_logic;
	-- signal N5_1_43 : std_logic;
	FA1509 : full_adder port map (N4_0_42,N4_1_42,N4_2_42,N5_0_42,N5_1_43);
-- In matrix 4 adding FA to column 42 
	-- signal N5_2_42 : std_logic;
	-- signal N5_3_43 : std_logic;
	FA1510 : full_adder port map (N4_3_42,N4_4_42,N4_5_42,N5_2_42,N5_3_43);
-- In matrix 4 adding FA to column 42 
	-- signal N5_4_42 : std_logic;
	-- signal N5_5_43 : std_logic;
	FA1511 : full_adder port map (N4_6_42,N4_7_42,N4_8_42,N5_4_42,N5_5_43);
-- In matrix 4 adding FA to column 42 
	-- signal N5_6_42 : std_logic;
	-- signal N5_7_43 : std_logic;
	FA1512 : full_adder port map (N4_9_42,N4_10_42,N4_11_42,N5_6_42,N5_7_43);
-- In matrix 4 adding FA to column 42 
	-- signal N5_8_42 : std_logic;
	-- signal N5_9_43 : std_logic;
	FA1513 : full_adder port map (N4_12_42,N4_13_42,N4_14_42,N5_8_42,N5_9_43);
-- In matrix 4 adding FA to column 43 
	-- signal N5_0_43 : std_logic;
	-- signal N5_1_44 : std_logic;
	FA1514 : full_adder port map (N4_0_43,N4_1_43,N4_2_43,N5_0_43,N5_1_44);
-- In matrix 4 adding FA to column 43 
	-- signal N5_2_43 : std_logic;
	-- signal N5_3_44 : std_logic;
	FA1515 : full_adder port map (N4_3_43,N4_4_43,N4_5_43,N5_2_43,N5_3_44);
-- In matrix 4 adding FA to column 43 
	-- signal N5_4_43 : std_logic;
	-- signal N5_5_44 : std_logic;
	FA1516 : full_adder port map (N4_6_43,N4_7_43,N4_8_43,N5_4_43,N5_5_44);
-- In matrix 4 adding FA to column 43 
	-- signal N5_6_43 : std_logic;
	-- signal N5_7_44 : std_logic;
	FA1517 : full_adder port map (N4_9_43,N4_10_43,N4_11_43,N5_6_43,N5_7_44);
-- In matrix 4 adding FA to column 43 
	-- signal N5_8_43 : std_logic;
	-- signal N5_9_44 : std_logic;
	FA1518 : full_adder port map (N4_12_43,N4_13_43,N4_14_43,N5_8_43,N5_9_44);
-- In matrix 4 adding FA to column 44 
	-- signal N5_0_44 : std_logic;
	-- signal N5_1_45 : std_logic;
	FA1519 : full_adder port map (N4_0_44,N4_1_44,N4_2_44,N5_0_44,N5_1_45);
-- In matrix 4 adding FA to column 44 
	-- signal N5_2_44 : std_logic;
	-- signal N5_3_45 : std_logic;
	FA1520 : full_adder port map (N4_3_44,N4_4_44,N4_5_44,N5_2_44,N5_3_45);
-- In matrix 4 adding FA to column 44 
	-- signal N5_4_44 : std_logic;
	-- signal N5_5_45 : std_logic;
	FA1521 : full_adder port map (N4_6_44,N4_7_44,N4_8_44,N5_4_44,N5_5_45);
-- In matrix 4 adding FA to column 44 
	-- signal N5_6_44 : std_logic;
	-- signal N5_7_45 : std_logic;
	FA1522 : full_adder port map (N4_9_44,N4_10_44,N4_11_44,N5_6_44,N5_7_45);
-- In matrix 4 adding FA to column 44 
	-- signal N5_8_44 : std_logic;
	-- signal N5_9_45 : std_logic;
	FA1523 : full_adder port map (N4_12_44,N4_13_44,N4_14_44,N5_8_44,N5_9_45);
-- In matrix 4 adding FA to column 45 
	-- signal N5_0_45 : std_logic;
	-- signal N5_1_46 : std_logic;
	FA1524 : full_adder port map (N4_0_45,N4_1_45,N4_2_45,N5_0_45,N5_1_46);
-- In matrix 4 adding FA to column 45 
	-- signal N5_2_45 : std_logic;
	-- signal N5_3_46 : std_logic;
	FA1525 : full_adder port map (N4_3_45,N4_4_45,N4_5_45,N5_2_45,N5_3_46);
-- In matrix 4 adding FA to column 45 
	-- signal N5_4_45 : std_logic;
	-- signal N5_5_46 : std_logic;
	FA1526 : full_adder port map (N4_6_45,N4_7_45,N4_8_45,N5_4_45,N5_5_46);
-- In matrix 4 adding FA to column 45 
	-- signal N5_6_45 : std_logic;
	-- signal N5_7_46 : std_logic;
	FA1527 : full_adder port map (N4_9_45,N4_10_45,N4_11_45,N5_6_45,N5_7_46);
-- In matrix 4 adding FA to column 45 
	-- signal N5_8_45 : std_logic;
	-- signal N5_9_46 : std_logic;
	FA1528 : full_adder port map (N4_12_45,N4_13_45,N4_14_45,N5_8_45,N5_9_46);
-- In matrix 4 adding FA to column 46 
	-- signal N5_0_46 : std_logic;
	-- signal N5_1_47 : std_logic;
	FA1529 : full_adder port map (N4_0_46,N4_1_46,N4_2_46,N5_0_46,N5_1_47);
-- In matrix 4 adding FA to column 46 
	-- signal N5_2_46 : std_logic;
	-- signal N5_3_47 : std_logic;
	FA1530 : full_adder port map (N4_3_46,N4_4_46,N4_5_46,N5_2_46,N5_3_47);
-- In matrix 4 adding FA to column 46 
	-- signal N5_4_46 : std_logic;
	-- signal N5_5_47 : std_logic;
	FA1531 : full_adder port map (N4_6_46,N4_7_46,N4_8_46,N5_4_46,N5_5_47);
-- In matrix 4 adding FA to column 46 
	-- signal N5_6_46 : std_logic;
	-- signal N5_7_47 : std_logic;
	FA1532 : full_adder port map (N4_9_46,N4_10_46,N4_11_46,N5_6_46,N5_7_47);
-- In matrix 4 adding FA to column 46 
	-- signal N5_8_46 : std_logic;
	-- signal N5_9_47 : std_logic;
	FA1533 : full_adder port map (N4_12_46,N4_13_46,N4_14_46,N5_8_46,N5_9_47);
-- In matrix 4 adding FA to column 47 
	-- signal N5_0_47 : std_logic;
	-- signal N5_1_48 : std_logic;
	FA1534 : full_adder port map (N4_0_47,N4_1_47,N4_2_47,N5_0_47,N5_1_48);
-- In matrix 4 adding FA to column 47 
	-- signal N5_2_47 : std_logic;
	-- signal N5_3_48 : std_logic;
	FA1535 : full_adder port map (N4_3_47,N4_4_47,N4_5_47,N5_2_47,N5_3_48);
-- In matrix 4 adding FA to column 47 
	-- signal N5_4_47 : std_logic;
	-- signal N5_5_48 : std_logic;
	FA1536 : full_adder port map (N4_6_47,N4_7_47,N4_8_47,N5_4_47,N5_5_48);
-- In matrix 4 adding FA to column 47 
	-- signal N5_6_47 : std_logic;
	-- signal N5_7_48 : std_logic;
	FA1537 : full_adder port map (N4_9_47,N4_10_47,N4_11_47,N5_6_47,N5_7_48);
-- In matrix 4 adding FA to column 47 
	-- signal N5_8_47 : std_logic;
	-- signal N5_9_48 : std_logic;
	FA1538 : full_adder port map (N4_12_47,N4_13_47,N4_14_47,N5_8_47,N5_9_48);
-- In matrix 4 adding FA to column 48 
	-- signal N5_0_48 : std_logic;
	-- signal N5_1_49 : std_logic;
	FA1539 : full_adder port map (N4_0_48,N4_1_48,N4_2_48,N5_0_48,N5_1_49);
-- In matrix 4 adding FA to column 48 
	-- signal N5_2_48 : std_logic;
	-- signal N5_3_49 : std_logic;
	FA1540 : full_adder port map (N4_3_48,N4_4_48,N4_5_48,N5_2_48,N5_3_49);
-- In matrix 4 adding FA to column 48 
	-- signal N5_4_48 : std_logic;
	-- signal N5_5_49 : std_logic;
	FA1541 : full_adder port map (N4_6_48,N4_7_48,N4_8_48,N5_4_48,N5_5_49);
-- In matrix 4 adding FA to column 48 
	-- signal N5_6_48 : std_logic;
	-- signal N5_7_49 : std_logic;
	FA1542 : full_adder port map (N4_9_48,N4_10_48,N4_11_48,N5_6_48,N5_7_49);
-- In matrix 4 adding FA to column 48 
	-- signal N5_8_48 : std_logic;
	-- signal N5_9_49 : std_logic;
	FA1543 : full_adder port map (N4_12_48,N4_13_48,N4_14_48,N5_8_48,N5_9_49);
-- In matrix 4 adding FA to column 49 
	-- signal N5_0_49 : std_logic;
	-- signal N5_1_50 : std_logic;
	FA1544 : full_adder port map (N4_0_49,N4_1_49,N4_2_49,N5_0_49,N5_1_50);
-- In matrix 4 adding FA to column 49 
	-- signal N5_2_49 : std_logic;
	-- signal N5_3_50 : std_logic;
	FA1545 : full_adder port map (N4_3_49,N4_4_49,N4_5_49,N5_2_49,N5_3_50);
-- In matrix 4 adding FA to column 49 
	-- signal N5_4_49 : std_logic;
	-- signal N5_5_50 : std_logic;
	FA1546 : full_adder port map (N4_6_49,N4_7_49,N4_8_49,N5_4_49,N5_5_50);
-- In matrix 4 adding FA to column 49 
	-- signal N5_6_49 : std_logic;
	-- signal N5_7_50 : std_logic;
	FA1547 : full_adder port map (N4_9_49,N4_10_49,N4_11_49,N5_6_49,N5_7_50);
-- In matrix 4 adding FA to column 49 
	-- signal N5_8_49 : std_logic;
	-- signal N5_9_50 : std_logic;
	FA1548 : full_adder port map (N4_12_49,N4_13_49,N4_14_49,N5_8_49,N5_9_50);
-- In matrix 4 adding FA to column 50 
	-- signal N5_0_50 : std_logic;
	-- signal N5_1_51 : std_logic;
	FA1549 : full_adder port map (N4_0_50,N4_1_50,N4_2_50,N5_0_50,N5_1_51);
-- In matrix 4 adding FA to column 50 
	-- signal N5_2_50 : std_logic;
	-- signal N5_3_51 : std_logic;
	FA1550 : full_adder port map (N4_3_50,N4_4_50,N4_5_50,N5_2_50,N5_3_51);
-- In matrix 4 adding FA to column 50 
	-- signal N5_4_50 : std_logic;
	-- signal N5_5_51 : std_logic;
	FA1551 : full_adder port map (N4_6_50,N4_7_50,N4_8_50,N5_4_50,N5_5_51);
-- In matrix 4 adding FA to column 50 
	-- signal N5_6_50 : std_logic;
	-- signal N5_7_51 : std_logic;
	FA1552 : full_adder port map (N4_9_50,N4_10_50,N4_11_50,N5_6_50,N5_7_51);
-- In matrix 4 adding FA to column 50 
	-- signal N5_8_50 : std_logic;
	-- signal N5_9_51 : std_logic;
	FA1553 : full_adder port map (N4_12_50,N4_13_50,N4_14_50,N5_8_50,N5_9_51);
-- In matrix 4 adding FA to column 51 
	-- signal N5_0_51 : std_logic;
	-- signal N5_1_52 : std_logic;
	FA1554 : full_adder port map (N4_0_51,N4_1_51,N4_2_51,N5_0_51,N5_1_52);
-- In matrix 4 adding FA to column 51 
	-- signal N5_2_51 : std_logic;
	-- signal N5_3_52 : std_logic;
	FA1555 : full_adder port map (N4_3_51,N4_4_51,N4_5_51,N5_2_51,N5_3_52);
-- In matrix 4 adding FA to column 51 
	-- signal N5_4_51 : std_logic;
	-- signal N5_5_52 : std_logic;
	FA1556 : full_adder port map (N4_6_51,N4_7_51,N4_8_51,N5_4_51,N5_5_52);
-- In matrix 4 adding FA to column 51 
	-- signal N5_6_51 : std_logic;
	-- signal N5_7_52 : std_logic;
	FA1557 : full_adder port map (N4_9_51,N4_10_51,N4_11_51,N5_6_51,N5_7_52);
-- In matrix 4 adding FA to column 51 
	-- signal N5_8_51 : std_logic;
	-- signal N5_9_52 : std_logic;
	FA1558 : full_adder port map (N4_12_51,N4_13_51,N4_14_51,N5_8_51,N5_9_52);
-- In matrix 4 adding FA to column 52 
	-- signal N5_0_52 : std_logic;
	-- signal N5_1_53 : std_logic;
	FA1559 : full_adder port map (N4_0_52,N4_1_52,N4_2_52,N5_0_52,N5_1_53);
-- In matrix 4 adding FA to column 52 
	-- signal N5_2_52 : std_logic;
	-- signal N5_3_53 : std_logic;
	FA1560 : full_adder port map (N4_3_52,N4_4_52,N4_5_52,N5_2_52,N5_3_53);
-- In matrix 4 adding FA to column 52 
	-- signal N5_4_52 : std_logic;
	-- signal N5_5_53 : std_logic;
	FA1561 : full_adder port map (N4_6_52,N4_7_52,N4_8_52,N5_4_52,N5_5_53);
-- In matrix 4 adding FA to column 52 
	-- signal N5_6_52 : std_logic;
	-- signal N5_7_53 : std_logic;
	FA1562 : full_adder port map (N4_9_52,N4_10_52,N4_11_52,N5_6_52,N5_7_53);
-- In matrix 4 adding FA to column 52 
	-- signal N5_8_52 : std_logic;
	-- signal N5_9_53 : std_logic;
	FA1563 : full_adder port map (N4_12_52,N4_13_52,N4_14_52,N5_8_52,N5_9_53);
-- In matrix 4 adding FA to column 53 
	-- signal N5_0_53 : std_logic;
	-- signal N5_1_54 : std_logic;
	FA1564 : full_adder port map (N4_0_53,N4_1_53,N4_2_53,N5_0_53,N5_1_54);
-- In matrix 4 adding FA to column 53 
	-- signal N5_2_53 : std_logic;
	-- signal N5_3_54 : std_logic;
	FA1565 : full_adder port map (N4_3_53,N4_4_53,N4_5_53,N5_2_53,N5_3_54);
-- In matrix 4 adding FA to column 53 
	-- signal N5_4_53 : std_logic;
	-- signal N5_5_54 : std_logic;
	FA1566 : full_adder port map (N4_6_53,N4_7_53,N4_8_53,N5_4_53,N5_5_54);
-- In matrix 4 adding FA to column 53 
	-- signal N5_6_53 : std_logic;
	-- signal N5_7_54 : std_logic;
	FA1567 : full_adder port map (N4_9_53,N4_10_53,N4_11_53,N5_6_53,N5_7_54);
-- In matrix 4 adding FA to column 53 
	-- signal N5_8_53 : std_logic;
	-- signal N5_9_54 : std_logic;
	FA1568 : full_adder port map (N4_12_53,N4_13_53,N4_14_53,N5_8_53,N5_9_54);
-- In matrix 4 adding FA to column 54 
	-- signal N5_0_54 : std_logic;
	-- signal N5_1_55 : std_logic;
	FA1569 : full_adder port map (N4_0_54,N4_1_54,N4_2_54,N5_0_54,N5_1_55);
-- In matrix 4 adding FA to column 54 
	-- signal N5_2_54 : std_logic;
	-- signal N5_3_55 : std_logic;
	FA1570 : full_adder port map (N4_3_54,N4_4_54,N4_5_54,N5_2_54,N5_3_55);
-- In matrix 4 adding FA to column 54 
	-- signal N5_4_54 : std_logic;
	-- signal N5_5_55 : std_logic;
	FA1571 : full_adder port map (N4_6_54,N4_7_54,N4_8_54,N5_4_54,N5_5_55);
-- In matrix 4 adding FA to column 54 
	-- signal N5_6_54 : std_logic;
	-- signal N5_7_55 : std_logic;
	FA1572 : full_adder port map (N4_9_54,N4_10_54,N4_11_54,N5_6_54,N5_7_55);
-- In matrix 4 adding FA to column 54 
	-- signal N5_8_54 : std_logic;
	-- signal N5_9_55 : std_logic;
	FA1573 : full_adder port map (N4_12_54,N4_13_54,N4_14_54,N5_8_54,N5_9_55);
-- In matrix 4 adding FA to column 55 
	-- signal N5_0_55 : std_logic;
	-- signal N5_1_56 : std_logic;
	FA1574 : full_adder port map (N4_0_55,N4_1_55,N4_2_55,N5_0_55,N5_1_56);
-- In matrix 4 adding FA to column 55 
	-- signal N5_2_55 : std_logic;
	-- signal N5_3_56 : std_logic;
	FA1575 : full_adder port map (N4_3_55,N4_4_55,N4_5_55,N5_2_55,N5_3_56);
-- In matrix 4 adding FA to column 55 
	-- signal N5_4_55 : std_logic;
	-- signal N5_5_56 : std_logic;
	FA1576 : full_adder port map (N4_6_55,N4_7_55,N4_8_55,N5_4_55,N5_5_56);
-- In matrix 4 adding FA to column 55 
	-- signal N5_6_55 : std_logic;
	-- signal N5_7_56 : std_logic;
	FA1577 : full_adder port map (N4_9_55,N4_10_55,N4_11_55,N5_6_55,N5_7_56);
-- In matrix 4 adding FA to column 55 
	-- signal N5_8_55 : std_logic;
	-- signal N5_9_56 : std_logic;
	FA1578 : full_adder port map (N4_12_55,N4_13_55,N4_14_55,N5_8_55,N5_9_56);
-- In matrix 4 adding FA to column 56 
	-- signal N5_0_56 : std_logic;
	-- signal N5_1_57 : std_logic;
	FA1579 : full_adder port map (N4_0_56,N4_1_56,N4_2_56,N5_0_56,N5_1_57);
-- In matrix 4 adding FA to column 56 
	-- signal N5_2_56 : std_logic;
	-- signal N5_3_57 : std_logic;
	FA1580 : full_adder port map (N4_3_56,N4_4_56,N4_5_56,N5_2_56,N5_3_57);
-- In matrix 4 adding FA to column 56 
	-- signal N5_4_56 : std_logic;
	-- signal N5_5_57 : std_logic;
	FA1581 : full_adder port map (N4_6_56,N4_7_56,N4_8_56,N5_4_56,N5_5_57);
-- In matrix 4 adding FA to column 56 
	-- signal N5_6_56 : std_logic;
	-- signal N5_7_57 : std_logic;
	FA1582 : full_adder port map (N4_9_56,N4_10_56,N4_11_56,N5_6_56,N5_7_57);
-- In matrix 4 adding FA to column 56 
	-- signal N5_8_56 : std_logic;
	-- signal N5_9_57 : std_logic;
	FA1583 : full_adder port map (N4_12_56,N4_13_56,N4_14_56,N5_8_56,N5_9_57);
-- In matrix 4 adding FA to column 57 
	-- signal N5_0_57 : std_logic;
	-- signal N5_1_58 : std_logic;
	FA1584 : full_adder port map (N4_0_57,N4_1_57,N4_2_57,N5_0_57,N5_1_58);
-- In matrix 4 adding FA to column 57 
	-- signal N5_2_57 : std_logic;
	-- signal N5_3_58 : std_logic;
	FA1585 : full_adder port map (N4_3_57,N4_4_57,N4_5_57,N5_2_57,N5_3_58);
-- In matrix 4 adding FA to column 57 
	-- signal N5_4_57 : std_logic;
	-- signal N5_5_58 : std_logic;
	FA1586 : full_adder port map (N4_6_57,N4_7_57,N4_8_57,N5_4_57,N5_5_58);
-- In matrix 4 adding FA to column 57 
	-- signal N5_6_57 : std_logic;
	-- signal N5_7_58 : std_logic;
	FA1587 : full_adder port map (N4_9_57,N4_10_57,N4_11_57,N5_6_57,N5_7_58);
-- In matrix 4 adding FA to column 57 
	-- signal N5_8_57 : std_logic;
	-- signal N5_9_58 : std_logic;
	FA1588 : full_adder port map (N4_12_57,N4_13_57,N4_14_57,N5_8_57,N5_9_58);
-- In matrix 4 adding FA to column 58 
	-- signal N5_0_58 : std_logic;
	-- signal N5_1_59 : std_logic;
	FA1589 : full_adder port map (N4_0_58,N4_1_58,N4_2_58,N5_0_58,N5_1_59);
-- In matrix 4 adding FA to column 58 
	-- signal N5_2_58 : std_logic;
	-- signal N5_3_59 : std_logic;
	FA1590 : full_adder port map (N4_3_58,N4_4_58,N4_5_58,N5_2_58,N5_3_59);
-- In matrix 4 adding FA to column 58 
	-- signal N5_4_58 : std_logic;
	-- signal N5_5_59 : std_logic;
	FA1591 : full_adder port map (N4_6_58,N4_7_58,N4_8_58,N5_4_58,N5_5_59);
-- In matrix 4 adding FA to column 58 
	-- signal N5_6_58 : std_logic;
	-- signal N5_7_59 : std_logic;
	FA1592 : full_adder port map (N4_9_58,N4_10_58,N4_11_58,N5_6_58,N5_7_59);
-- In matrix 4 adding FA to column 58 
	-- signal N5_8_58 : std_logic;
	-- signal N5_9_59 : std_logic;
	FA1593 : full_adder port map (N4_12_58,N4_13_58,N4_14_58,N5_8_58,N5_9_59);
-- In matrix 4 adding FA to column 59 
	-- signal N5_0_59 : std_logic;
	-- signal N5_1_60 : std_logic;
	FA1594 : full_adder port map (N4_0_59,N4_1_59,N4_2_59,N5_0_59,N5_1_60);
-- In matrix 4 adding FA to column 59 
	-- signal N5_2_59 : std_logic;
	-- signal N5_3_60 : std_logic;
	FA1595 : full_adder port map (N4_3_59,N4_4_59,N4_5_59,N5_2_59,N5_3_60);
-- In matrix 4 adding FA to column 59 
	-- signal N5_4_59 : std_logic;
	-- signal N5_5_60 : std_logic;
	FA1596 : full_adder port map (N4_6_59,N4_7_59,N4_8_59,N5_4_59,N5_5_60);
-- In matrix 4 adding FA to column 59 
	-- signal N5_6_59 : std_logic;
	-- signal N5_7_60 : std_logic;
	FA1597 : full_adder port map (N4_9_59,N4_10_59,N4_11_59,N5_6_59,N5_7_60);
-- In matrix 4 adding FA to column 59 
	-- signal N5_8_59 : std_logic;
	-- signal N5_9_60 : std_logic;
	FA1598 : full_adder port map (N4_12_59,N4_13_59,N4_14_59,N5_8_59,N5_9_60);
-- In matrix 4 adding FA to column 60 
	-- signal N5_0_60 : std_logic;
	-- signal N5_1_61 : std_logic;
	FA1599 : full_adder port map (N4_0_60,N4_1_60,N4_2_60,N5_0_60,N5_1_61);
-- In matrix 4 adding FA to column 60 
	-- signal N5_2_60 : std_logic;
	-- signal N5_3_61 : std_logic;
	FA1600 : full_adder port map (N4_3_60,N4_4_60,N4_5_60,N5_2_60,N5_3_61);
-- In matrix 4 adding FA to column 60 
	-- signal N5_4_60 : std_logic;
	-- signal N5_5_61 : std_logic;
	FA1601 : full_adder port map (N4_6_60,N4_7_60,N4_8_60,N5_4_60,N5_5_61);
-- In matrix 4 adding FA to column 60 
	-- signal N5_6_60 : std_logic;
	-- signal N5_7_61 : std_logic;
	FA1602 : full_adder port map (N4_9_60,N4_10_60,N4_11_60,N5_6_60,N5_7_61);
-- In matrix 4 adding FA to column 60 
	-- signal N5_8_60 : std_logic;
	-- signal N5_9_61 : std_logic;
	FA1603 : full_adder port map (N4_12_60,N4_13_60,N4_14_60,N5_8_60,N5_9_61);
-- In matrix 4 adding FA to column 61 
	-- signal N5_0_61 : std_logic;
	-- signal N5_1_62 : std_logic;
	FA1604 : full_adder port map (N4_0_61,N4_1_61,N4_2_61,N5_0_61,N5_1_62);
-- In matrix 4 adding FA to column 61 
	-- signal N5_2_61 : std_logic;
	-- signal N5_3_62 : std_logic;
	FA1605 : full_adder port map (N4_3_61,N4_4_61,N4_5_61,N5_2_61,N5_3_62);
-- In matrix 4 adding FA to column 61 
	-- signal N5_4_61 : std_logic;
	-- signal N5_5_62 : std_logic;
	FA1606 : full_adder port map (N4_6_61,N4_7_61,N4_8_61,N5_4_61,N5_5_62);
-- In matrix 4 adding FA to column 61 
	-- signal N5_6_61 : std_logic;
	-- signal N5_7_62 : std_logic;
	FA1607 : full_adder port map (N4_9_61,N4_10_61,N4_11_61,N5_6_61,N5_7_62);
-- In matrix 4 adding FA to column 61 
	-- signal N5_8_61 : std_logic;
	-- signal N5_9_62 : std_logic;
	FA1608 : full_adder port map (N4_12_61,N4_13_61,N4_14_61,N5_8_61,N5_9_62);
-- In matrix 4 adding FA to column 62 
	-- signal N5_0_62 : std_logic;
	-- signal N5_1_63 : std_logic;
	FA1609 : full_adder port map (N4_0_62,N4_1_62,N4_2_62,N5_0_62,N5_1_63);
-- In matrix 4 adding FA to column 62 
	-- signal N5_2_62 : std_logic;
	-- signal N5_3_63 : std_logic;
	FA1610 : full_adder port map (N4_3_62,N4_4_62,N4_5_62,N5_2_62,N5_3_63);
-- In matrix 4 adding FA to column 62 
	-- signal N5_4_62 : std_logic;
	-- signal N5_5_63 : std_logic;
	FA1611 : full_adder port map (N4_6_62,N4_7_62,N4_8_62,N5_4_62,N5_5_63);
-- In matrix 4 adding FA to column 62 
	-- signal N5_6_62 : std_logic;
	-- signal N5_7_63 : std_logic;
	FA1612 : full_adder port map (N4_9_62,N4_10_62,N4_11_62,N5_6_62,N5_7_63);
-- In matrix 4 adding FA to column 62 
	-- signal N5_8_62 : std_logic;
	-- signal N5_9_63 : std_logic;
	FA1613 : full_adder port map (N4_12_62,N4_13_62,N4_14_62,N5_8_62,N5_9_63);
-- In matrix 4 adding FA to column 63 
	-- signal N5_0_63 : std_logic;
	-- signal N5_1_64 : std_logic;
	FA1614 : full_adder port map (N4_0_63,N4_1_63,N4_2_63,N5_0_63,N5_1_64);
-- In matrix 4 adding FA to column 63 
	-- signal N5_2_63 : std_logic;
	-- signal N5_3_64 : std_logic;
	FA1615 : full_adder port map (N4_3_63,N4_4_63,N4_5_63,N5_2_63,N5_3_64);
-- In matrix 4 adding FA to column 63 
	-- signal N5_4_63 : std_logic;
	-- signal N5_5_64 : std_logic;
	FA1616 : full_adder port map (N4_6_63,N4_7_63,N4_8_63,N5_4_63,N5_5_64);
-- In matrix 4 adding FA to column 63 
	-- signal N5_6_63 : std_logic;
	-- signal N5_7_64 : std_logic;
	FA1617 : full_adder port map (N4_9_63,N4_10_63,N4_11_63,N5_6_63,N5_7_64);
-- In matrix 4 adding FA to column 63 
	-- signal N5_8_63 : std_logic;
	-- signal N5_9_64 : std_logic;
	FA1618 : full_adder port map (N4_12_63,N4_13_63,N4_14_63,N5_8_63,N5_9_64);
-- In matrix 4 adding FA to column 64 
	-- signal N5_0_64 : std_logic;
	-- signal N5_1_65 : std_logic;
	FA1619 : full_adder port map (N4_0_64,N4_1_64,N4_2_64,N5_0_64,N5_1_65);
-- In matrix 4 adding FA to column 64 
	-- signal N5_2_64 : std_logic;
	-- signal N5_3_65 : std_logic;
	FA1620 : full_adder port map (N4_3_64,N4_4_64,N4_5_64,N5_2_64,N5_3_65);
-- In matrix 4 adding FA to column 64 
	-- signal N5_4_64 : std_logic;
	-- signal N5_5_65 : std_logic;
	FA1621 : full_adder port map (N4_6_64,N4_7_64,N4_8_64,N5_4_64,N5_5_65);
-- In matrix 4 adding FA to column 64 
	-- signal N5_6_64 : std_logic;
	-- signal N5_7_65 : std_logic;
	FA1622 : full_adder port map (N4_9_64,N4_10_64,N4_11_64,N5_6_64,N5_7_65);
-- In matrix 4 adding FA to column 64 
	-- signal N5_8_64 : std_logic;
	-- signal N5_9_65 : std_logic;
	FA1623 : full_adder port map (N4_12_64,N4_13_64,N4_14_64,N5_8_64,N5_9_65);
-- In matrix 4 adding FA to column 65 
	-- signal N5_0_65 : std_logic;
	-- signal N5_1_66 : std_logic;
	FA1624 : full_adder port map (N4_0_65,N4_1_65,N4_2_65,N5_0_65,N5_1_66);
-- In matrix 4 adding FA to column 65 
	-- signal N5_2_65 : std_logic;
	-- signal N5_3_66 : std_logic;
	FA1625 : full_adder port map (N4_3_65,N4_4_65,N4_5_65,N5_2_65,N5_3_66);
-- In matrix 4 adding FA to column 65 
	-- signal N5_4_65 : std_logic;
	-- signal N5_5_66 : std_logic;
	FA1626 : full_adder port map (N4_6_65,N4_7_65,N4_8_65,N5_4_65,N5_5_66);
-- In matrix 4 adding FA to column 65 
	-- signal N5_6_65 : std_logic;
	-- signal N5_7_66 : std_logic;
	FA1627 : full_adder port map (N4_9_65,N4_10_65,N4_11_65,N5_6_65,N5_7_66);
-- In matrix 4 adding FA to column 65 
	-- signal N5_8_65 : std_logic;
	-- signal N5_9_66 : std_logic;
	FA1628 : full_adder port map (N4_12_65,N4_13_65,N4_14_65,N5_8_65,N5_9_66);
-- In matrix 4 adding FA to column 66 
	-- signal N5_0_66 : std_logic;
	-- signal N5_1_67 : std_logic;
	FA1629 : full_adder port map (N4_0_66,N4_1_66,N4_2_66,N5_0_66,N5_1_67);
-- In matrix 4 adding FA to column 66 
	-- signal N5_2_66 : std_logic;
	-- signal N5_3_67 : std_logic;
	FA1630 : full_adder port map (N4_3_66,N4_4_66,N4_5_66,N5_2_66,N5_3_67);
-- In matrix 4 adding FA to column 66 
	-- signal N5_4_66 : std_logic;
	-- signal N5_5_67 : std_logic;
	FA1631 : full_adder port map (N4_6_66,N4_7_66,N4_8_66,N5_4_66,N5_5_67);
-- In matrix 4 adding FA to column 66 
	-- signal N5_6_66 : std_logic;
	-- signal N5_7_67 : std_logic;
	FA1632 : full_adder port map (N4_9_66,N4_10_66,N4_11_66,N5_6_66,N5_7_67);
-- In matrix 4 adding FA to column 66 
	-- signal N5_8_66 : std_logic;
	-- signal N5_9_67 : std_logic;
	FA1633 : full_adder port map (N4_12_66,N4_13_66,N4_14_66,N5_8_66,N5_9_67);
-- In matrix 4 adding FA to column 67 
	-- signal N5_0_67 : std_logic;
	-- signal N5_1_68 : std_logic;
	FA1634 : full_adder port map (N4_0_67,N4_1_67,N4_2_67,N5_0_67,N5_1_68);
-- In matrix 4 adding FA to column 67 
	-- signal N5_2_67 : std_logic;
	-- signal N5_3_68 : std_logic;
	FA1635 : full_adder port map (N4_3_67,N4_4_67,N4_5_67,N5_2_67,N5_3_68);
-- In matrix 4 adding FA to column 67 
	-- signal N5_4_67 : std_logic;
	-- signal N5_5_68 : std_logic;
	FA1636 : full_adder port map (N4_6_67,N4_7_67,N4_8_67,N5_4_67,N5_5_68);
-- In matrix 4 adding FA to column 67 
	-- signal N5_6_67 : std_logic;
	-- signal N5_7_68 : std_logic;
	FA1637 : full_adder port map (N4_9_67,N4_10_67,N4_11_67,N5_6_67,N5_7_68);
-- In matrix 4 adding FA to column 67 
	-- signal N5_8_67 : std_logic;
	-- signal N5_9_68 : std_logic;
	FA1638 : full_adder port map (N4_12_67,N4_13_67,N4_14_67,N5_8_67,N5_9_68);
-- In matrix 4 adding FA to column 68 
	-- signal N5_0_68 : std_logic;
	-- signal N5_1_69 : std_logic;
	FA1639 : full_adder port map (N4_0_68,N4_1_68,N4_2_68,N5_0_68,N5_1_69);
-- In matrix 4 adding FA to column 68 
	-- signal N5_2_68 : std_logic;
	-- signal N5_3_69 : std_logic;
	FA1640 : full_adder port map (N4_3_68,N4_4_68,N4_5_68,N5_2_68,N5_3_69);
-- In matrix 4 adding FA to column 68 
	-- signal N5_4_68 : std_logic;
	-- signal N5_5_69 : std_logic;
	FA1641 : full_adder port map (N4_6_68,N4_7_68,N4_8_68,N5_4_68,N5_5_69);
-- In matrix 4 adding FA to column 68 
	-- signal N5_6_68 : std_logic;
	-- signal N5_7_69 : std_logic;
	FA1642 : full_adder port map (N4_9_68,N4_10_68,N4_11_68,N5_6_68,N5_7_69);
-- In matrix 4 adding FA to column 68 
	-- signal N5_8_68 : std_logic;
	-- signal N5_9_69 : std_logic;
	FA1643 : full_adder port map (N4_12_68,N4_13_68,N4_14_68,N5_8_68,N5_9_69);
-- In matrix 4 adding FA to column 69 
	-- signal N5_0_69 : std_logic;
	-- signal N5_1_70 : std_logic;
	FA1644 : full_adder port map (N4_0_69,N4_1_69,N4_2_69,N5_0_69,N5_1_70);
-- In matrix 4 adding FA to column 69 
	-- signal N5_2_69 : std_logic;
	-- signal N5_3_70 : std_logic;
	FA1645 : full_adder port map (N4_3_69,N4_4_69,N4_5_69,N5_2_69,N5_3_70);
-- In matrix 4 adding FA to column 69 
	-- signal N5_4_69 : std_logic;
	-- signal N5_5_70 : std_logic;
	FA1646 : full_adder port map (N4_6_69,N4_7_69,N4_8_69,N5_4_69,N5_5_70);
-- In matrix 4 adding FA to column 69 
	-- signal N5_6_69 : std_logic;
	-- signal N5_7_70 : std_logic;
	FA1647 : full_adder port map (N4_9_69,N4_10_69,N4_11_69,N5_6_69,N5_7_70);
-- In matrix 4 adding FA to column 69 
	-- signal N5_8_69 : std_logic;
	-- signal N5_9_70 : std_logic;
	FA1648 : full_adder port map (N4_12_69,N4_13_69,N4_14_69,N5_8_69,N5_9_70);
-- In matrix 4 adding FA to column 70 
	-- signal N5_0_70 : std_logic;
	-- signal N5_1_71 : std_logic;
	FA1649 : full_adder port map (N4_0_70,N4_1_70,N4_2_70,N5_0_70,N5_1_71);
-- In matrix 4 adding FA to column 70 
	-- signal N5_2_70 : std_logic;
	-- signal N5_3_71 : std_logic;
	FA1650 : full_adder port map (N4_3_70,N4_4_70,N4_5_70,N5_2_70,N5_3_71);
-- In matrix 4 adding FA to column 70 
	-- signal N5_4_70 : std_logic;
	-- signal N5_5_71 : std_logic;
	FA1651 : full_adder port map (N4_6_70,N4_7_70,N4_8_70,N5_4_70,N5_5_71);
-- In matrix 4 adding FA to column 70 
	-- signal N5_6_70 : std_logic;
	-- signal N5_7_71 : std_logic;
	FA1652 : full_adder port map (N4_9_70,N4_10_70,N4_11_70,N5_6_70,N5_7_71);
-- In matrix 4 adding FA to column 70 
	-- signal N5_8_70 : std_logic;
	-- signal N5_9_71 : std_logic;
	FA1653 : full_adder port map (N4_12_70,N4_13_70,N4_14_70,N5_8_70,N5_9_71);
-- In matrix 4 adding FA to column 71 
	-- signal N5_0_71 : std_logic;
	-- signal N5_1_72 : std_logic;
	FA1654 : full_adder port map (N4_0_71,N4_1_71,N4_2_71,N5_0_71,N5_1_72);
-- In matrix 4 adding FA to column 71 
	-- signal N5_2_71 : std_logic;
	-- signal N5_3_72 : std_logic;
	FA1655 : full_adder port map (N4_3_71,N4_4_71,N4_5_71,N5_2_71,N5_3_72);
-- In matrix 4 adding FA to column 71 
	-- signal N5_4_71 : std_logic;
	-- signal N5_5_72 : std_logic;
	FA1656 : full_adder port map (N4_6_71,N4_7_71,N4_8_71,N5_4_71,N5_5_72);
-- In matrix 4 adding FA to column 71 
	-- signal N5_6_71 : std_logic;
	-- signal N5_7_72 : std_logic;
	FA1657 : full_adder port map (N4_9_71,N4_10_71,N4_11_71,N5_6_71,N5_7_72);
-- In matrix 4 adding FA to column 71 
	-- signal N5_8_71 : std_logic;
	-- signal N5_9_72 : std_logic;
	FA1658 : full_adder port map (N4_12_71,N4_13_71,N4_14_71,N5_8_71,N5_9_72);
-- In matrix 4 adding FA to column 72 
	-- signal N5_0_72 : std_logic;
	-- signal N5_1_73 : std_logic;
	FA1659 : full_adder port map (N4_0_72,N4_1_72,N4_2_72,N5_0_72,N5_1_73);
-- In matrix 4 adding FA to column 72 
	-- signal N5_2_72 : std_logic;
	-- signal N5_3_73 : std_logic;
	FA1660 : full_adder port map (N4_3_72,N4_4_72,N4_5_72,N5_2_72,N5_3_73);
-- In matrix 4 adding FA to column 72 
	-- signal N5_4_72 : std_logic;
	-- signal N5_5_73 : std_logic;
	FA1661 : full_adder port map (N4_6_72,N4_7_72,N4_8_72,N5_4_72,N5_5_73);
-- In matrix 4 adding FA to column 72 
	-- signal N5_6_72 : std_logic;
	-- signal N5_7_73 : std_logic;
	FA1662 : full_adder port map (N4_9_72,N4_10_72,N4_11_72,N5_6_72,N5_7_73);
-- In matrix 4 adding FA to column 72 
	-- signal N5_8_72 : std_logic;
	-- signal N5_9_73 : std_logic;
	FA1663 : full_adder port map (N4_12_72,N4_13_72,N4_14_72,N5_8_72,N5_9_73);
-- In matrix 4 adding FA to column 73 
	-- signal N5_0_73 : std_logic;
	-- signal N5_1_74 : std_logic;
	FA1664 : full_adder port map (N4_0_73,N4_1_73,N4_2_73,N5_0_73,N5_1_74);
-- In matrix 4 adding FA to column 73 
	-- signal N5_2_73 : std_logic;
	-- signal N5_3_74 : std_logic;
	FA1665 : full_adder port map (N4_3_73,N4_4_73,N4_5_73,N5_2_73,N5_3_74);
-- In matrix 4 adding FA to column 73 
	-- signal N5_4_73 : std_logic;
	-- signal N5_5_74 : std_logic;
	FA1666 : full_adder port map (N4_6_73,N4_7_73,N4_8_73,N5_4_73,N5_5_74);
-- In matrix 4 adding FA to column 73 
	-- signal N5_6_73 : std_logic;
	-- signal N5_7_74 : std_logic;
	FA1667 : full_adder port map (N4_9_73,N4_10_73,N4_11_73,N5_6_73,N5_7_74);
-- In matrix 4 adding FA to column 73 
	-- signal N5_8_73 : std_logic;
	-- signal N5_9_74 : std_logic;
	FA1668 : full_adder port map (N4_12_73,N4_13_73,N4_14_73,N5_8_73,N5_9_74);
-- In matrix 4 adding FA to column 74 
	-- signal N5_0_74 : std_logic;
	-- signal N5_1_75 : std_logic;
	FA1669 : full_adder port map (N4_0_74,N4_1_74,N4_2_74,N5_0_74,N5_1_75);
-- In matrix 4 adding FA to column 74 
	-- signal N5_2_74 : std_logic;
	-- signal N5_3_75 : std_logic;
	FA1670 : full_adder port map (N4_3_74,N4_4_74,N4_5_74,N5_2_74,N5_3_75);
-- In matrix 4 adding FA to column 74 
	-- signal N5_4_74 : std_logic;
	-- signal N5_5_75 : std_logic;
	FA1671 : full_adder port map (N4_6_74,N4_7_74,N4_8_74,N5_4_74,N5_5_75);
-- In matrix 4 adding FA to column 74 
	-- signal N5_6_74 : std_logic;
	-- signal N5_7_75 : std_logic;
	FA1672 : full_adder port map (N4_9_74,N4_10_74,N4_11_74,N5_6_74,N5_7_75);
-- In matrix 4 adding FA to column 74 
	-- signal N5_8_74 : std_logic;
	-- signal N5_9_75 : std_logic;
	FA1673 : full_adder port map (N4_12_74,N4_13_74,N4_14_74,N5_8_74,N5_9_75);
-- In matrix 4 adding FA to column 75 
	-- signal N5_0_75 : std_logic;
	-- signal N5_1_76 : std_logic;
	FA1674 : full_adder port map (N4_0_75,N4_1_75,N4_2_75,N5_0_75,N5_1_76);
-- In matrix 4 adding FA to column 75 
	-- signal N5_2_75 : std_logic;
	-- signal N5_3_76 : std_logic;
	FA1675 : full_adder port map (N4_3_75,N4_4_75,N4_5_75,N5_2_75,N5_3_76);
-- In matrix 4 adding FA to column 75 
	-- signal N5_4_75 : std_logic;
	-- signal N5_5_76 : std_logic;
	FA1676 : full_adder port map (N4_6_75,N4_7_75,N4_8_75,N5_4_75,N5_5_76);
-- In matrix 4 adding FA to column 75 
	-- signal N5_6_75 : std_logic;
	-- signal N5_7_76 : std_logic;
	FA1677 : full_adder port map (N4_9_75,N4_10_75,N4_11_75,N5_6_75,N5_7_76);
-- In matrix 4 adding FA to column 75 
	-- signal N5_8_75 : std_logic;
	-- signal N5_9_76 : std_logic;
	FA1678 : full_adder port map (N4_12_75,N4_13_75,N4_14_75,N5_8_75,N5_9_76);
-- In matrix 4 adding FA to column 76 
	-- signal N5_0_76 : std_logic;
	-- signal N5_1_77 : std_logic;
	FA1679 : full_adder port map (N4_0_76,N4_1_76,N4_2_76,N5_0_76,N5_1_77);
-- In matrix 4 adding FA to column 76 
	-- signal N5_2_76 : std_logic;
	-- signal N5_3_77 : std_logic;
	FA1680 : full_adder port map (N4_3_76,N4_4_76,N4_5_76,N5_2_76,N5_3_77);
-- In matrix 4 adding FA to column 76 
	-- signal N5_4_76 : std_logic;
	-- signal N5_5_77 : std_logic;
	FA1681 : full_adder port map (N4_6_76,N4_7_76,N4_8_76,N5_4_76,N5_5_77);
-- In matrix 4 adding FA to column 76 
	-- signal N5_6_76 : std_logic;
	-- signal N5_7_77 : std_logic;
	FA1682 : full_adder port map (N4_9_76,N4_10_76,N4_11_76,N5_6_76,N5_7_77);
-- In matrix 4 adding FA to column 76 
	-- signal N5_8_76 : std_logic;
	-- signal N5_9_77 : std_logic;
	FA1683 : full_adder port map (N4_12_76,N4_13_76,N4_14_76,N5_8_76,N5_9_77);
-- In matrix 4 adding FA to column 77 
	-- signal N5_0_77 : std_logic;
	-- signal N5_1_78 : std_logic;
	FA1684 : full_adder port map (N4_0_77,N4_1_77,N4_2_77,N5_0_77,N5_1_78);
-- In matrix 4 adding FA to column 77 
	-- signal N5_2_77 : std_logic;
	-- signal N5_3_78 : std_logic;
	FA1685 : full_adder port map (N4_3_77,N4_4_77,N4_5_77,N5_2_77,N5_3_78);
-- In matrix 4 adding FA to column 77 
	-- signal N5_4_77 : std_logic;
	-- signal N5_5_78 : std_logic;
	FA1686 : full_adder port map (N4_6_77,N4_7_77,N4_8_77,N5_4_77,N5_5_78);
-- In matrix 4 adding FA to column 77 
	-- signal N5_6_77 : std_logic;
	-- signal N5_7_78 : std_logic;
	FA1687 : full_adder port map (N4_9_77,N4_10_77,N4_11_77,N5_6_77,N5_7_78);
-- In matrix 4 adding FA to column 77 
	-- signal N5_8_77 : std_logic;
	-- signal N5_9_78 : std_logic;
	FA1688 : full_adder port map (N4_12_77,N4_13_77,N4_14_77,N5_8_77,N5_9_78);
-- In matrix 4 adding FA to column 78 
	-- signal N5_0_78 : std_logic;
	-- signal N5_1_79 : std_logic;
	FA1689 : full_adder port map (N4_0_78,N4_1_78,N4_2_78,N5_0_78,N5_1_79);
-- In matrix 4 adding FA to column 78 
	-- signal N5_2_78 : std_logic;
	-- signal N5_3_79 : std_logic;
	FA1690 : full_adder port map (N4_3_78,N4_4_78,N4_5_78,N5_2_78,N5_3_79);
-- In matrix 4 adding FA to column 78 
	-- signal N5_4_78 : std_logic;
	-- signal N5_5_79 : std_logic;
	FA1691 : full_adder port map (N4_6_78,N4_7_78,N4_8_78,N5_4_78,N5_5_79);
-- In matrix 4 adding FA to column 78 
	-- signal N5_6_78 : std_logic;
	-- signal N5_7_79 : std_logic;
	FA1692 : full_adder port map (N4_9_78,N4_10_78,N4_11_78,N5_6_78,N5_7_79);
-- In matrix 4 adding FA to column 78 
	-- signal N5_8_78 : std_logic;
	-- signal N5_9_79 : std_logic;
	FA1693 : full_adder port map (N4_12_78,N4_13_78,N4_14_78,N5_8_78,N5_9_79);
-- In matrix 4 adding FA to column 79 
	-- signal N5_0_79 : std_logic;
	-- signal N5_1_80 : std_logic;
	FA1694 : full_adder port map (N4_0_79,N4_1_79,N4_2_79,N5_0_79,N5_1_80);
-- In matrix 4 adding FA to column 79 
	-- signal N5_2_79 : std_logic;
	-- signal N5_3_80 : std_logic;
	FA1695 : full_adder port map (N4_3_79,N4_4_79,N4_5_79,N5_2_79,N5_3_80);
-- In matrix 4 adding FA to column 79 
	-- signal N5_4_79 : std_logic;
	-- signal N5_5_80 : std_logic;
	FA1696 : full_adder port map (N4_6_79,N4_7_79,N4_8_79,N5_4_79,N5_5_80);
-- In matrix 4 adding FA to column 79 
	-- signal N5_6_79 : std_logic;
	-- signal N5_7_80 : std_logic;
	FA1697 : full_adder port map (N4_9_79,N4_10_79,N4_11_79,N5_6_79,N5_7_80);
-- In matrix 4 adding FA to column 79 
	-- signal N5_8_79 : std_logic;
	-- signal N5_9_80 : std_logic;
	FA1698 : full_adder port map (N4_12_79,N4_13_79,N4_14_79,N5_8_79,N5_9_80);
-- In matrix 4 adding FA to column 80 
	-- signal N5_0_80 : std_logic;
	-- signal N5_1_81 : std_logic;
	FA1699 : full_adder port map (N4_0_80,N4_1_80,N4_2_80,N5_0_80,N5_1_81);
-- In matrix 4 adding FA to column 80 
	-- signal N5_2_80 : std_logic;
	-- signal N5_3_81 : std_logic;
	FA1700 : full_adder port map (N4_3_80,N4_4_80,N4_5_80,N5_2_80,N5_3_81);
-- In matrix 4 adding FA to column 80 
	-- signal N5_4_80 : std_logic;
	-- signal N5_5_81 : std_logic;
	FA1701 : full_adder port map (N4_6_80,N4_7_80,N4_8_80,N5_4_80,N5_5_81);
-- In matrix 4 adding FA to column 80 
	-- signal N5_6_80 : std_logic;
	-- signal N5_7_81 : std_logic;
	FA1702 : full_adder port map (N4_9_80,N4_10_80,N4_11_80,N5_6_80,N5_7_81);
-- In matrix 4 adding FA to column 80 
	-- signal N5_8_80 : std_logic;
	-- signal N5_9_81 : std_logic;
	FA1703 : full_adder port map (N4_12_80,N4_13_80,N4_14_80,N5_8_80,N5_9_81);
-- In matrix 4 adding FA to column 81 
	-- signal N5_0_81 : std_logic;
	-- signal N5_1_82 : std_logic;
	FA1704 : full_adder port map (N4_0_81,N4_1_81,N4_2_81,N5_0_81,N5_1_82);
-- In matrix 4 adding FA to column 81 
	-- signal N5_2_81 : std_logic;
	-- signal N5_3_82 : std_logic;
	FA1705 : full_adder port map (N4_3_81,N4_4_81,N4_5_81,N5_2_81,N5_3_82);
-- In matrix 4 adding FA to column 81 
	-- signal N5_4_81 : std_logic;
	-- signal N5_5_82 : std_logic;
	FA1706 : full_adder port map (N4_6_81,N4_7_81,N4_8_81,N5_4_81,N5_5_82);
-- In matrix 4 adding FA to column 81 
	-- signal N5_6_81 : std_logic;
	-- signal N5_7_82 : std_logic;
	FA1707 : full_adder port map (N4_9_81,N4_10_81,N4_11_81,N5_6_81,N5_7_82);
-- In matrix 4 adding FA to column 81 
	-- signal N5_8_81 : std_logic;
	-- signal N5_9_82 : std_logic;
	FA1708 : full_adder port map (N4_12_81,N4_13_81,N4_14_81,N5_8_81,N5_9_82);
-- In matrix 4 adding FA to column 82 
	-- signal N5_0_82 : std_logic;
	-- signal N5_1_83 : std_logic;
	FA1709 : full_adder port map (N4_0_82,N4_1_82,N4_2_82,N5_0_82,N5_1_83);
-- In matrix 4 adding FA to column 82 
	-- signal N5_2_82 : std_logic;
	-- signal N5_3_83 : std_logic;
	FA1710 : full_adder port map (N4_3_82,N4_4_82,N4_5_82,N5_2_82,N5_3_83);
-- In matrix 4 adding FA to column 82 
	-- signal N5_4_82 : std_logic;
	-- signal N5_5_83 : std_logic;
	FA1711 : full_adder port map (N4_6_82,N4_7_82,N4_8_82,N5_4_82,N5_5_83);
-- In matrix 4 adding FA to column 82 
	-- signal N5_6_82 : std_logic;
	-- signal N5_7_83 : std_logic;
	FA1712 : full_adder port map (N4_9_82,N4_10_82,N4_11_82,N5_6_82,N5_7_83);
-- In matrix 4 adding FA to column 82 
	-- signal N5_8_82 : std_logic;
	-- signal N5_9_83 : std_logic;
	FA1713 : full_adder port map (N4_12_82,N4_13_82,N4_14_82,N5_8_82,N5_9_83);
-- In matrix 4 adding FA to column 83 
	-- signal N5_0_83 : std_logic;
	-- signal N5_1_84 : std_logic;
	FA1714 : full_adder port map (N0_52_83,N4_0_83,N4_1_83,N5_0_83,N5_1_84);
-- In matrix 4 adding FA to column 83 
	-- signal N5_2_83 : std_logic;
	-- signal N5_3_84 : std_logic;
	FA1715 : full_adder port map (N4_2_83,N4_3_83,N4_4_83,N5_2_83,N5_3_84);
-- In matrix 4 adding FA to column 83 
	-- signal N5_4_83 : std_logic;
	-- signal N5_5_84 : std_logic;
	FA1716 : full_adder port map (N4_5_83,N4_6_83,N4_7_83,N5_4_83,N5_5_84);
-- In matrix 4 adding FA to column 83 
	-- signal N5_6_83 : std_logic;
	-- signal N5_7_84 : std_logic;
	FA1717 : full_adder port map (N4_8_83,N4_9_83,N4_10_83,N5_6_83,N5_7_84);
-- In matrix 4 adding FA to column 83 
	-- signal N5_8_83 : std_logic;
	-- signal N5_9_84 : std_logic;
	FA1718 : full_adder port map (N4_11_83,N4_12_83,N4_13_83,N5_8_83,N5_9_84);
-- In matrix 4 adding FA to column 84 
	-- signal N5_0_84 : std_logic;
	-- signal N5_1_85 : std_logic;
	FA1719 : full_adder port map (N0_50_84,N0_51_84,N0_52_84,N5_0_84,N5_1_85);
-- In matrix 4 adding FA to column 84 
	-- signal N5_2_84 : std_logic;
	-- signal N5_3_85 : std_logic;
	FA1720 : full_adder port map (N4_0_84,N4_1_84,N4_2_84,N5_2_84,N5_3_85);
-- In matrix 4 adding FA to column 84 
	-- signal N5_4_84 : std_logic;
	-- signal N5_5_85 : std_logic;
	FA1721 : full_adder port map (N4_3_84,N4_4_84,N4_5_84,N5_4_84,N5_5_85);
-- In matrix 4 adding FA to column 84 
	-- signal N5_6_84 : std_logic;
	-- signal N5_7_85 : std_logic;
	FA1722 : full_adder port map (N4_6_84,N4_7_84,N4_8_84,N5_6_84,N5_7_85);
-- In matrix 4 adding FA to column 84 
	-- signal N5_8_84 : std_logic;
	-- signal N5_9_85 : std_logic;
	FA1723 : full_adder port map (N4_9_84,N4_10_84,N4_11_84,N5_8_84,N5_9_85);
-- In matrix 4 adding FA to column 85 
	-- signal N5_0_85 : std_logic;
	-- signal N5_1_86 : std_logic;
	FA1724 : full_adder port map (N0_48_85,N0_49_85,N0_50_85,N5_0_85,N5_1_86);
-- In matrix 4 adding FA to column 85 
	-- signal N5_2_85 : std_logic;
	-- signal N5_3_86 : std_logic;
	FA1725 : full_adder port map (N0_51_85,N0_52_85,N4_0_85,N5_2_85,N5_3_86);
-- In matrix 4 adding FA to column 85 
	-- signal N5_4_85 : std_logic;
	-- signal N5_5_86 : std_logic;
	FA1726 : full_adder port map (N4_1_85,N4_2_85,N4_3_85,N5_4_85,N5_5_86);
-- In matrix 4 adding FA to column 85 
	-- signal N5_6_85 : std_logic;
	-- signal N5_7_86 : std_logic;
	FA1727 : full_adder port map (N4_4_85,N4_5_85,N4_6_85,N5_6_85,N5_7_86);
-- In matrix 4 adding FA to column 85 
	-- signal N5_8_85 : std_logic;
	-- signal N5_9_86 : std_logic;
	FA1728 : full_adder port map (N4_7_85,N4_8_85,N4_9_85,N5_8_85,N5_9_86);
-- In matrix 4 adding FA to column 86 
	-- signal N5_0_86 : std_logic;
	-- signal N5_1_87 : std_logic;
	FA1729 : full_adder port map (N0_46_86,N0_47_86,N0_48_86,N5_0_86,N5_1_87);
-- In matrix 4 adding FA to column 86 
	-- signal N5_2_86 : std_logic;
	-- signal N5_3_87 : std_logic;
	FA1730 : full_adder port map (N0_49_86,N0_50_86,N0_51_86,N5_2_86,N5_3_87);
-- In matrix 4 adding FA to column 86 
	-- signal N5_4_86 : std_logic;
	-- signal N5_5_87 : std_logic;
	FA1731 : full_adder port map (N0_52_86,N4_0_86,N4_1_86,N5_4_86,N5_5_87);
-- In matrix 4 adding FA to column 86 
	-- signal N5_6_86 : std_logic;
	-- signal N5_7_87 : std_logic;
	FA1732 : full_adder port map (N4_2_86,N4_3_86,N4_4_86,N5_6_86,N5_7_87);
-- In matrix 4 adding FA to column 86 
	-- signal N5_8_86 : std_logic;
	-- signal N5_9_87 : std_logic;
	FA1733 : full_adder port map (N4_5_86,N4_6_86,N4_7_86,N5_8_86,N5_9_87);
-- In matrix 4 adding FA to column 87 
	-- signal N5_0_87 : std_logic;
	-- signal N5_1_88 : std_logic;
	FA1734 : full_adder port map (N0_44_87,N0_45_87,N0_46_87,N5_0_87,N5_1_88);
-- In matrix 4 adding FA to column 87 
	-- signal N5_2_87 : std_logic;
	-- signal N5_3_88 : std_logic;
	FA1735 : full_adder port map (N0_47_87,N0_48_87,N0_49_87,N5_2_87,N5_3_88);
-- In matrix 4 adding FA to column 87 
	-- signal N5_4_87 : std_logic;
	-- signal N5_5_88 : std_logic;
	FA1736 : full_adder port map (N0_50_87,N0_51_87,N0_52_87,N5_4_87,N5_5_88);
-- In matrix 4 adding FA to column 87 
	-- signal N5_6_87 : std_logic;
	-- signal N5_7_88 : std_logic;
	FA1737 : full_adder port map (N4_0_87,N4_1_87,N4_2_87,N5_6_87,N5_7_88);
-- In matrix 4 adding FA to column 87 
	-- signal N5_8_87 : std_logic;
	-- signal N5_9_88 : std_logic;
	FA1738 : full_adder port map (N4_3_87,N4_4_87,N4_5_87,N5_8_87,N5_9_88);
-- In matrix 4 adding FA to column 88 
	-- signal N5_0_88 : std_logic;
	-- signal N5_1_89 : std_logic;
	FA1739 : full_adder port map (N0_42_88,N0_43_88,N0_44_88,N5_0_88,N5_1_89);
-- In matrix 4 adding FA to column 88 
	-- signal N5_2_88 : std_logic;
	-- signal N5_3_89 : std_logic;
	FA1740 : full_adder port map (N0_45_88,N0_46_88,N0_47_88,N5_2_88,N5_3_89);
-- In matrix 4 adding FA to column 88 
	-- signal N5_4_88 : std_logic;
	-- signal N5_5_89 : std_logic;
	FA1741 : full_adder port map (N0_48_88,N0_49_88,N0_50_88,N5_4_88,N5_5_89);
-- In matrix 4 adding FA to column 88 
	-- signal N5_6_88 : std_logic;
	-- signal N5_7_89 : std_logic;
	FA1742 : full_adder port map (N0_51_88,N0_52_88,N4_0_88,N5_6_88,N5_7_89);
-- In matrix 4 adding FA to column 88 
	-- signal N5_8_88 : std_logic;
	-- signal N5_9_89 : std_logic;
	FA1743 : full_adder port map (N4_1_88,N4_2_88,N4_3_88,N5_8_88,N5_9_89);
-- In matrix 4 adding FA to column 89 
	-- signal N5_0_89 : std_logic;
	-- signal N5_1_90 : std_logic;
	FA1744 : full_adder port map (N0_40_89,N0_41_89,N0_42_89,N5_0_89,N5_1_90);
-- In matrix 4 adding FA to column 89 
	-- signal N5_2_89 : std_logic;
	-- signal N5_3_90 : std_logic;
	FA1745 : full_adder port map (N0_43_89,N0_44_89,N0_45_89,N5_2_89,N5_3_90);
-- In matrix 4 adding FA to column 89 
	-- signal N5_4_89 : std_logic;
	-- signal N5_5_90 : std_logic;
	FA1746 : full_adder port map (N0_46_89,N0_47_89,N0_48_89,N5_4_89,N5_5_90);
-- In matrix 4 adding FA to column 89 
	-- signal N5_6_89 : std_logic;
	-- signal N5_7_90 : std_logic;
	FA1747 : full_adder port map (N0_49_89,N0_50_89,N0_51_89,N5_6_89,N5_7_90);
-- In matrix 4 adding FA to column 89 
	-- signal N5_8_89 : std_logic;
	-- signal N5_9_90 : std_logic;
	FA1748 : full_adder port map (N0_52_89,N4_0_89,N4_1_89,N5_8_89,N5_9_90);
-- In matrix 4 adding FA to column 90 
	-- signal N5_0_90 : std_logic;
	-- signal N5_1_91 : std_logic;
	FA1749 : full_adder port map (N0_38_90,N0_39_90,N0_40_90,N5_0_90,N5_1_91);
-- In matrix 4 adding FA to column 90 
	-- signal N5_2_90 : std_logic;
	-- signal N5_3_91 : std_logic;
	FA1750 : full_adder port map (N0_41_90,N0_42_90,N0_43_90,N5_2_90,N5_3_91);
-- In matrix 4 adding FA to column 90 
	-- signal N5_4_90 : std_logic;
	-- signal N5_5_91 : std_logic;
	FA1751 : full_adder port map (N0_44_90,N0_45_90,N0_46_90,N5_4_90,N5_5_91);
-- In matrix 4 adding FA to column 90 
	-- signal N5_6_90 : std_logic;
	-- signal N5_7_91 : std_logic;
	FA1752 : full_adder port map (N0_47_90,N0_48_90,N0_49_90,N5_6_90,N5_7_91);
-- In matrix 4 adding FA to column 90 
	-- signal N5_8_90 : std_logic;
	-- signal N5_9_91 : std_logic;
	FA1753 : full_adder port map (N0_50_90,N0_51_90,N0_52_90,N5_8_90,N5_9_91);
-- In matrix 4 adding FA to column 91 
	-- signal N5_0_91 : std_logic;
	-- signal N5_1_92 : std_logic;
	FA1754 : full_adder port map (N0_39_91,N0_40_91,N0_41_91,N5_0_91,N5_1_92);
-- In matrix 4 adding FA to column 91 
	-- signal N5_2_91 : std_logic;
	-- signal N5_3_92 : std_logic;
	FA1755 : full_adder port map (N0_42_91,N0_43_91,N0_44_91,N5_2_91,N5_3_92);
-- In matrix 4 adding FA to column 91 
	-- signal N5_4_91 : std_logic;
	-- signal N5_5_92 : std_logic;
	FA1756 : full_adder port map (N0_45_91,N0_46_91,N0_47_91,N5_4_91,N5_5_92);
-- In matrix 4 adding FA to column 91 
	-- signal N5_6_91 : std_logic;
	-- signal N5_7_92 : std_logic;
	FA1757 : full_adder port map (N0_48_91,N0_49_91,N0_50_91,N5_6_91,N5_7_92);
-- In matrix 4 adding FA to column 92 
	-- signal N5_0_92 : std_logic;
	-- signal N5_1_93 : std_logic;
	FA1758 : full_adder port map (N0_40_92,N0_41_92,N0_42_92,N5_0_92,N5_1_93);
-- In matrix 4 adding FA to column 92 
	-- signal N5_2_92 : std_logic;
	-- signal N5_3_93 : std_logic;
	FA1759 : full_adder port map (N0_43_92,N0_44_92,N0_45_92,N5_2_92,N5_3_93);
-- In matrix 4 adding FA to column 92 
	-- signal N5_4_92 : std_logic;
	-- signal N5_5_93 : std_logic;
	FA1760 : full_adder port map (N0_46_92,N0_47_92,N0_48_92,N5_4_92,N5_5_93);
-- In matrix 4 adding FA to column 93 
	-- signal N5_0_93 : std_logic;
	-- signal N5_1_94 : std_logic;
	FA1761 : full_adder port map (N0_41_93,N0_42_93,N0_43_93,N5_0_93,N5_1_94);
-- In matrix 4 adding FA to column 93 
	-- signal N5_2_93 : std_logic;
	-- signal N5_3_94 : std_logic;
	FA1762 : full_adder port map (N0_44_93,N0_45_93,N0_46_93,N5_2_93,N5_3_94);
-- In matrix 4 adding FA to column 94 
	-- signal N5_0_94 : std_logic;
	-- signal N5_1_95 : std_logic;
	FA1763 : full_adder port map (N0_42_94,N0_43_94,N0_44_94,N5_0_94,N5_1_95);
	-- Elements from matrix 5 
-- In matrix 5 adding HA to column 8 
	-- signal N6_0_8 : std_logic;
	-- signal N6_1_9 : std_logic;
	HA44 : half_adder port map (N0_0_8,N0_1_8,N6_0_8,N6_1_9);
-- In matrix 5 adding FA to column 9 
	-- signal N6_0_9 : std_logic;
	-- signal N6_1_10 : std_logic;
	FA1764 : full_adder port map (N0_0_9,N0_1_9,N0_2_9,N6_0_9,N6_1_10);
-- In matrix 5 adding HA to column 9 
	-- signal N6_2_9 : std_logic;
	-- signal N6_3_10 : std_logic;
	HA45 : half_adder port map (N0_3_9,N0_4_9,N6_2_9,N6_3_10);
-- In matrix 5 adding FA to column 10 
	-- signal N6_0_10 : std_logic;
	-- signal N6_1_11 : std_logic;
	FA1765 : full_adder port map (N0_0_10,N0_1_10,N0_2_10,N6_0_10,N6_1_11);
-- In matrix 5 adding FA to column 10 
	-- signal N6_2_10 : std_logic;
	-- signal N6_3_11 : std_logic;
	FA1766 : full_adder port map (N0_3_10,N0_4_10,N0_5_10,N6_2_10,N6_3_11);
-- In matrix 5 adding HA to column 10 
	-- signal N6_4_10 : std_logic;
	-- signal N6_5_11 : std_logic;
	HA46 : half_adder port map (N0_6_10,N0_7_10,N6_4_10,N6_5_11);
-- In matrix 5 adding FA to column 11 
	-- signal N6_0_11 : std_logic;
	-- signal N6_1_12 : std_logic;
	FA1767 : full_adder port map (N0_2_11,N0_3_11,N0_4_11,N6_0_11,N6_1_12);
-- In matrix 5 adding FA to column 11 
	-- signal N6_2_11 : std_logic;
	-- signal N6_3_12 : std_logic;
	FA1768 : full_adder port map (N0_5_11,N0_6_11,N0_7_11,N6_2_11,N6_3_12);
-- In matrix 5 adding FA to column 11 
	-- signal N6_4_11 : std_logic;
	-- signal N6_5_12 : std_logic;
	FA1769 : full_adder port map (N0_8_11,N0_9_11,N0_10_11,N6_4_11,N6_5_12);
-- In matrix 5 adding FA to column 12 
	-- signal N6_0_12 : std_logic;
	-- signal N6_1_13 : std_logic;
	FA1770 : full_adder port map (N0_5_12,N0_6_12,N0_7_12,N6_0_12,N6_1_13);
-- In matrix 5 adding FA to column 12 
	-- signal N6_2_12 : std_logic;
	-- signal N6_3_13 : std_logic;
	FA1771 : full_adder port map (N0_8_12,N0_9_12,N0_10_12,N6_2_12,N6_3_13);
-- In matrix 5 adding FA to column 12 
	-- signal N6_4_12 : std_logic;
	-- signal N6_5_13 : std_logic;
	FA1772 : full_adder port map (N0_11_12,N0_12_12,N5_0_12,N6_4_12,N6_5_13);
-- In matrix 5 adding FA to column 13 
	-- signal N6_0_13 : std_logic;
	-- signal N6_1_14 : std_logic;
	FA1773 : full_adder port map (N0_8_13,N0_9_13,N0_10_13,N6_0_13,N6_1_14);
-- In matrix 5 adding FA to column 13 
	-- signal N6_2_13 : std_logic;
	-- signal N6_3_14 : std_logic;
	FA1774 : full_adder port map (N0_11_13,N0_12_13,N0_13_13,N6_2_13,N6_3_14);
-- In matrix 5 adding FA to column 13 
	-- signal N6_4_13 : std_logic;
	-- signal N6_5_14 : std_logic;
	FA1775 : full_adder port map (N5_0_13,N5_1_13,N5_2_13,N6_4_13,N6_5_14);
-- In matrix 5 adding FA to column 14 
	-- signal N6_0_14 : std_logic;
	-- signal N6_1_15 : std_logic;
	FA1776 : full_adder port map (N0_11_14,N0_12_14,N0_13_14,N6_0_14,N6_1_15);
-- In matrix 5 adding FA to column 14 
	-- signal N6_2_14 : std_logic;
	-- signal N6_3_15 : std_logic;
	FA1777 : full_adder port map (N0_14_14,N5_0_14,N5_1_14,N6_2_14,N6_3_15);
-- In matrix 5 adding FA to column 14 
	-- signal N6_4_14 : std_logic;
	-- signal N6_5_15 : std_logic;
	FA1778 : full_adder port map (N5_2_14,N5_3_14,N5_4_14,N6_4_14,N6_5_15);
-- In matrix 5 adding FA to column 15 
	-- signal N6_0_15 : std_logic;
	-- signal N6_1_16 : std_logic;
	FA1779 : full_adder port map (N0_14_15,N0_15_15,N5_0_15,N6_0_15,N6_1_16);
-- In matrix 5 adding FA to column 15 
	-- signal N6_2_15 : std_logic;
	-- signal N6_3_16 : std_logic;
	FA1780 : full_adder port map (N5_1_15,N5_2_15,N5_3_15,N6_2_15,N6_3_16);
-- In matrix 5 adding FA to column 15 
	-- signal N6_4_15 : std_logic;
	-- signal N6_5_16 : std_logic;
	FA1781 : full_adder port map (N5_4_15,N5_5_15,N5_6_15,N6_4_15,N6_5_16);
-- In matrix 5 adding FA to column 16 
	-- signal N6_0_16 : std_logic;
	-- signal N6_1_17 : std_logic;
	FA1782 : full_adder port map (N4_0_16,N5_0_16,N5_1_16,N6_0_16,N6_1_17);
-- In matrix 5 adding FA to column 16 
	-- signal N6_2_16 : std_logic;
	-- signal N6_3_17 : std_logic;
	FA1783 : full_adder port map (N5_2_16,N5_3_16,N5_4_16,N6_2_16,N6_3_17);
-- In matrix 5 adding FA to column 16 
	-- signal N6_4_16 : std_logic;
	-- signal N6_5_17 : std_logic;
	FA1784 : full_adder port map (N5_5_16,N5_6_16,N5_7_16,N6_4_16,N6_5_17);
-- In matrix 5 adding FA to column 17 
	-- signal N6_0_17 : std_logic;
	-- signal N6_1_18 : std_logic;
	FA1785 : full_adder port map (N4_2_17,N5_0_17,N5_1_17,N6_0_17,N6_1_18);
-- In matrix 5 adding FA to column 17 
	-- signal N6_2_17 : std_logic;
	-- signal N6_3_18 : std_logic;
	FA1786 : full_adder port map (N5_2_17,N5_3_17,N5_4_17,N6_2_17,N6_3_18);
-- In matrix 5 adding FA to column 17 
	-- signal N6_4_17 : std_logic;
	-- signal N6_5_18 : std_logic;
	FA1787 : full_adder port map (N5_5_17,N5_6_17,N5_7_17,N6_4_17,N6_5_18);
-- In matrix 5 adding FA to column 18 
	-- signal N6_0_18 : std_logic;
	-- signal N6_1_19 : std_logic;
	FA1788 : full_adder port map (N4_4_18,N5_0_18,N5_1_18,N6_0_18,N6_1_19);
-- In matrix 5 adding FA to column 18 
	-- signal N6_2_18 : std_logic;
	-- signal N6_3_19 : std_logic;
	FA1789 : full_adder port map (N5_2_18,N5_3_18,N5_4_18,N6_2_18,N6_3_19);
-- In matrix 5 adding FA to column 18 
	-- signal N6_4_18 : std_logic;
	-- signal N6_5_19 : std_logic;
	FA1790 : full_adder port map (N5_5_18,N5_6_18,N5_7_18,N6_4_18,N6_5_19);
-- In matrix 5 adding FA to column 19 
	-- signal N6_0_19 : std_logic;
	-- signal N6_1_20 : std_logic;
	FA1791 : full_adder port map (N4_6_19,N5_0_19,N5_1_19,N6_0_19,N6_1_20);
-- In matrix 5 adding FA to column 19 
	-- signal N6_2_19 : std_logic;
	-- signal N6_3_20 : std_logic;
	FA1792 : full_adder port map (N5_2_19,N5_3_19,N5_4_19,N6_2_19,N6_3_20);
-- In matrix 5 adding FA to column 19 
	-- signal N6_4_19 : std_logic;
	-- signal N6_5_20 : std_logic;
	FA1793 : full_adder port map (N5_5_19,N5_6_19,N5_7_19,N6_4_19,N6_5_20);
-- In matrix 5 adding FA to column 20 
	-- signal N6_0_20 : std_logic;
	-- signal N6_1_21 : std_logic;
	FA1794 : full_adder port map (N4_8_20,N5_0_20,N5_1_20,N6_0_20,N6_1_21);
-- In matrix 5 adding FA to column 20 
	-- signal N6_2_20 : std_logic;
	-- signal N6_3_21 : std_logic;
	FA1795 : full_adder port map (N5_2_20,N5_3_20,N5_4_20,N6_2_20,N6_3_21);
-- In matrix 5 adding FA to column 20 
	-- signal N6_4_20 : std_logic;
	-- signal N6_5_21 : std_logic;
	FA1796 : full_adder port map (N5_5_20,N5_6_20,N5_7_20,N6_4_20,N6_5_21);
-- In matrix 5 adding FA to column 21 
	-- signal N6_0_21 : std_logic;
	-- signal N6_1_22 : std_logic;
	FA1797 : full_adder port map (N4_10_21,N5_0_21,N5_1_21,N6_0_21,N6_1_22);
-- In matrix 5 adding FA to column 21 
	-- signal N6_2_21 : std_logic;
	-- signal N6_3_22 : std_logic;
	FA1798 : full_adder port map (N5_2_21,N5_3_21,N5_4_21,N6_2_21,N6_3_22);
-- In matrix 5 adding FA to column 21 
	-- signal N6_4_21 : std_logic;
	-- signal N6_5_22 : std_logic;
	FA1799 : full_adder port map (N5_5_21,N5_6_21,N5_7_21,N6_4_21,N6_5_22);
-- In matrix 5 adding FA to column 22 
	-- signal N6_0_22 : std_logic;
	-- signal N6_1_23 : std_logic;
	FA1800 : full_adder port map (N4_12_22,N5_0_22,N5_1_22,N6_0_22,N6_1_23);
-- In matrix 5 adding FA to column 22 
	-- signal N6_2_22 : std_logic;
	-- signal N6_3_23 : std_logic;
	FA1801 : full_adder port map (N5_2_22,N5_3_22,N5_4_22,N6_2_22,N6_3_23);
-- In matrix 5 adding FA to column 22 
	-- signal N6_4_22 : std_logic;
	-- signal N6_5_23 : std_logic;
	FA1802 : full_adder port map (N5_5_22,N5_6_22,N5_7_22,N6_4_22,N6_5_23);
-- In matrix 5 adding FA to column 23 
	-- signal N6_0_23 : std_logic;
	-- signal N6_1_24 : std_logic;
	FA1803 : full_adder port map (N4_14_23,N5_0_23,N5_1_23,N6_0_23,N6_1_24);
-- In matrix 5 adding FA to column 23 
	-- signal N6_2_23 : std_logic;
	-- signal N6_3_24 : std_logic;
	FA1804 : full_adder port map (N5_2_23,N5_3_23,N5_4_23,N6_2_23,N6_3_24);
-- In matrix 5 adding FA to column 23 
	-- signal N6_4_23 : std_logic;
	-- signal N6_5_24 : std_logic;
	FA1805 : full_adder port map (N5_5_23,N5_6_23,N5_7_23,N6_4_23,N6_5_24);
-- In matrix 5 adding FA to column 24 
	-- signal N6_0_24 : std_logic;
	-- signal N6_1_25 : std_logic;
	FA1806 : full_adder port map (N4_15_24,N5_0_24,N5_1_24,N6_0_24,N6_1_25);
-- In matrix 5 adding FA to column 24 
	-- signal N6_2_24 : std_logic;
	-- signal N6_3_25 : std_logic;
	FA1807 : full_adder port map (N5_2_24,N5_3_24,N5_4_24,N6_2_24,N6_3_25);
-- In matrix 5 adding FA to column 24 
	-- signal N6_4_24 : std_logic;
	-- signal N6_5_25 : std_logic;
	FA1808 : full_adder port map (N5_5_24,N5_6_24,N5_7_24,N6_4_24,N6_5_25);
-- In matrix 5 adding FA to column 25 
	-- signal N6_0_25 : std_logic;
	-- signal N6_1_26 : std_logic;
	FA1809 : full_adder port map (N4_15_25,N5_0_25,N5_1_25,N6_0_25,N6_1_26);
-- In matrix 5 adding FA to column 25 
	-- signal N6_2_25 : std_logic;
	-- signal N6_3_26 : std_logic;
	FA1810 : full_adder port map (N5_2_25,N5_3_25,N5_4_25,N6_2_25,N6_3_26);
-- In matrix 5 adding FA to column 25 
	-- signal N6_4_25 : std_logic;
	-- signal N6_5_26 : std_logic;
	FA1811 : full_adder port map (N5_5_25,N5_6_25,N5_7_25,N6_4_25,N6_5_26);
-- In matrix 5 adding FA to column 26 
	-- signal N6_0_26 : std_logic;
	-- signal N6_1_27 : std_logic;
	FA1812 : full_adder port map (N4_15_26,N5_0_26,N5_1_26,N6_0_26,N6_1_27);
-- In matrix 5 adding FA to column 26 
	-- signal N6_2_26 : std_logic;
	-- signal N6_3_27 : std_logic;
	FA1813 : full_adder port map (N5_2_26,N5_3_26,N5_4_26,N6_2_26,N6_3_27);
-- In matrix 5 adding FA to column 26 
	-- signal N6_4_26 : std_logic;
	-- signal N6_5_27 : std_logic;
	FA1814 : full_adder port map (N5_5_26,N5_6_26,N5_7_26,N6_4_26,N6_5_27);
-- In matrix 5 adding FA to column 27 
	-- signal N6_0_27 : std_logic;
	-- signal N6_1_28 : std_logic;
	FA1815 : full_adder port map (N4_15_27,N5_0_27,N5_1_27,N6_0_27,N6_1_28);
-- In matrix 5 adding FA to column 27 
	-- signal N6_2_27 : std_logic;
	-- signal N6_3_28 : std_logic;
	FA1816 : full_adder port map (N5_2_27,N5_3_27,N5_4_27,N6_2_27,N6_3_28);
-- In matrix 5 adding FA to column 27 
	-- signal N6_4_27 : std_logic;
	-- signal N6_5_28 : std_logic;
	FA1817 : full_adder port map (N5_5_27,N5_6_27,N5_7_27,N6_4_27,N6_5_28);
-- In matrix 5 adding FA to column 28 
	-- signal N6_0_28 : std_logic;
	-- signal N6_1_29 : std_logic;
	FA1818 : full_adder port map (N4_15_28,N5_0_28,N5_1_28,N6_0_28,N6_1_29);
-- In matrix 5 adding FA to column 28 
	-- signal N6_2_28 : std_logic;
	-- signal N6_3_29 : std_logic;
	FA1819 : full_adder port map (N5_2_28,N5_3_28,N5_4_28,N6_2_28,N6_3_29);
-- In matrix 5 adding FA to column 28 
	-- signal N6_4_28 : std_logic;
	-- signal N6_5_29 : std_logic;
	FA1820 : full_adder port map (N5_5_28,N5_6_28,N5_7_28,N6_4_28,N6_5_29);
-- In matrix 5 adding FA to column 29 
	-- signal N6_0_29 : std_logic;
	-- signal N6_1_30 : std_logic;
	FA1821 : full_adder port map (N4_15_29,N5_0_29,N5_1_29,N6_0_29,N6_1_30);
-- In matrix 5 adding FA to column 29 
	-- signal N6_2_29 : std_logic;
	-- signal N6_3_30 : std_logic;
	FA1822 : full_adder port map (N5_2_29,N5_3_29,N5_4_29,N6_2_29,N6_3_30);
-- In matrix 5 adding FA to column 29 
	-- signal N6_4_29 : std_logic;
	-- signal N6_5_30 : std_logic;
	FA1823 : full_adder port map (N5_5_29,N5_6_29,N5_7_29,N6_4_29,N6_5_30);
-- In matrix 5 adding FA to column 30 
	-- signal N6_0_30 : std_logic;
	-- signal N6_1_31 : std_logic;
	FA1824 : full_adder port map (N4_15_30,N5_0_30,N5_1_30,N6_0_30,N6_1_31);
-- In matrix 5 adding FA to column 30 
	-- signal N6_2_30 : std_logic;
	-- signal N6_3_31 : std_logic;
	FA1825 : full_adder port map (N5_2_30,N5_3_30,N5_4_30,N6_2_30,N6_3_31);
-- In matrix 5 adding FA to column 30 
	-- signal N6_4_30 : std_logic;
	-- signal N6_5_31 : std_logic;
	FA1826 : full_adder port map (N5_5_30,N5_6_30,N5_7_30,N6_4_30,N6_5_31);
-- In matrix 5 adding FA to column 31 
	-- signal N6_0_31 : std_logic;
	-- signal N6_1_32 : std_logic;
	FA1827 : full_adder port map (N4_15_31,N5_0_31,N5_1_31,N6_0_31,N6_1_32);
-- In matrix 5 adding FA to column 31 
	-- signal N6_2_31 : std_logic;
	-- signal N6_3_32 : std_logic;
	FA1828 : full_adder port map (N5_2_31,N5_3_31,N5_4_31,N6_2_31,N6_3_32);
-- In matrix 5 adding FA to column 31 
	-- signal N6_4_31 : std_logic;
	-- signal N6_5_32 : std_logic;
	FA1829 : full_adder port map (N5_5_31,N5_6_31,N5_7_31,N6_4_31,N6_5_32);
-- In matrix 5 adding FA to column 32 
	-- signal N6_0_32 : std_logic;
	-- signal N6_1_33 : std_logic;
	FA1830 : full_adder port map (N4_15_32,N5_0_32,N5_1_32,N6_0_32,N6_1_33);
-- In matrix 5 adding FA to column 32 
	-- signal N6_2_32 : std_logic;
	-- signal N6_3_33 : std_logic;
	FA1831 : full_adder port map (N5_2_32,N5_3_32,N5_4_32,N6_2_32,N6_3_33);
-- In matrix 5 adding FA to column 32 
	-- signal N6_4_32 : std_logic;
	-- signal N6_5_33 : std_logic;
	FA1832 : full_adder port map (N5_5_32,N5_6_32,N5_7_32,N6_4_32,N6_5_33);
-- In matrix 5 adding FA to column 33 
	-- signal N6_0_33 : std_logic;
	-- signal N6_1_34 : std_logic;
	FA1833 : full_adder port map (N4_15_33,N5_0_33,N5_1_33,N6_0_33,N6_1_34);
-- In matrix 5 adding FA to column 33 
	-- signal N6_2_33 : std_logic;
	-- signal N6_3_34 : std_logic;
	FA1834 : full_adder port map (N5_2_33,N5_3_33,N5_4_33,N6_2_33,N6_3_34);
-- In matrix 5 adding FA to column 33 
	-- signal N6_4_33 : std_logic;
	-- signal N6_5_34 : std_logic;
	FA1835 : full_adder port map (N5_5_33,N5_6_33,N5_7_33,N6_4_33,N6_5_34);
-- In matrix 5 adding FA to column 34 
	-- signal N6_0_34 : std_logic;
	-- signal N6_1_35 : std_logic;
	FA1836 : full_adder port map (N4_15_34,N5_0_34,N5_1_34,N6_0_34,N6_1_35);
-- In matrix 5 adding FA to column 34 
	-- signal N6_2_34 : std_logic;
	-- signal N6_3_35 : std_logic;
	FA1837 : full_adder port map (N5_2_34,N5_3_34,N5_4_34,N6_2_34,N6_3_35);
-- In matrix 5 adding FA to column 34 
	-- signal N6_4_34 : std_logic;
	-- signal N6_5_35 : std_logic;
	FA1838 : full_adder port map (N5_5_34,N5_6_34,N5_7_34,N6_4_34,N6_5_35);
-- In matrix 5 adding FA to column 35 
	-- signal N6_0_35 : std_logic;
	-- signal N6_1_36 : std_logic;
	FA1839 : full_adder port map (N4_15_35,N5_0_35,N5_1_35,N6_0_35,N6_1_36);
-- In matrix 5 adding FA to column 35 
	-- signal N6_2_35 : std_logic;
	-- signal N6_3_36 : std_logic;
	FA1840 : full_adder port map (N5_2_35,N5_3_35,N5_4_35,N6_2_35,N6_3_36);
-- In matrix 5 adding FA to column 35 
	-- signal N6_4_35 : std_logic;
	-- signal N6_5_36 : std_logic;
	FA1841 : full_adder port map (N5_5_35,N5_6_35,N5_7_35,N6_4_35,N6_5_36);
-- In matrix 5 adding FA to column 36 
	-- signal N6_0_36 : std_logic;
	-- signal N6_1_37 : std_logic;
	FA1842 : full_adder port map (N4_15_36,N5_0_36,N5_1_36,N6_0_36,N6_1_37);
-- In matrix 5 adding FA to column 36 
	-- signal N6_2_36 : std_logic;
	-- signal N6_3_37 : std_logic;
	FA1843 : full_adder port map (N5_2_36,N5_3_36,N5_4_36,N6_2_36,N6_3_37);
-- In matrix 5 adding FA to column 36 
	-- signal N6_4_36 : std_logic;
	-- signal N6_5_37 : std_logic;
	FA1844 : full_adder port map (N5_5_36,N5_6_36,N5_7_36,N6_4_36,N6_5_37);
-- In matrix 5 adding FA to column 37 
	-- signal N6_0_37 : std_logic;
	-- signal N6_1_38 : std_logic;
	FA1845 : full_adder port map (N4_15_37,N5_0_37,N5_1_37,N6_0_37,N6_1_38);
-- In matrix 5 adding FA to column 37 
	-- signal N6_2_37 : std_logic;
	-- signal N6_3_38 : std_logic;
	FA1846 : full_adder port map (N5_2_37,N5_3_37,N5_4_37,N6_2_37,N6_3_38);
-- In matrix 5 adding FA to column 37 
	-- signal N6_4_37 : std_logic;
	-- signal N6_5_38 : std_logic;
	FA1847 : full_adder port map (N5_5_37,N5_6_37,N5_7_37,N6_4_37,N6_5_38);
-- In matrix 5 adding FA to column 38 
	-- signal N6_0_38 : std_logic;
	-- signal N6_1_39 : std_logic;
	FA1848 : full_adder port map (N4_15_38,N5_0_38,N5_1_38,N6_0_38,N6_1_39);
-- In matrix 5 adding FA to column 38 
	-- signal N6_2_38 : std_logic;
	-- signal N6_3_39 : std_logic;
	FA1849 : full_adder port map (N5_2_38,N5_3_38,N5_4_38,N6_2_38,N6_3_39);
-- In matrix 5 adding FA to column 38 
	-- signal N6_4_38 : std_logic;
	-- signal N6_5_39 : std_logic;
	FA1850 : full_adder port map (N5_5_38,N5_6_38,N5_7_38,N6_4_38,N6_5_39);
-- In matrix 5 adding FA to column 39 
	-- signal N6_0_39 : std_logic;
	-- signal N6_1_40 : std_logic;
	FA1851 : full_adder port map (N4_15_39,N5_0_39,N5_1_39,N6_0_39,N6_1_40);
-- In matrix 5 adding FA to column 39 
	-- signal N6_2_39 : std_logic;
	-- signal N6_3_40 : std_logic;
	FA1852 : full_adder port map (N5_2_39,N5_3_39,N5_4_39,N6_2_39,N6_3_40);
-- In matrix 5 adding FA to column 39 
	-- signal N6_4_39 : std_logic;
	-- signal N6_5_40 : std_logic;
	FA1853 : full_adder port map (N5_5_39,N5_6_39,N5_7_39,N6_4_39,N6_5_40);
-- In matrix 5 adding FA to column 40 
	-- signal N6_0_40 : std_logic;
	-- signal N6_1_41 : std_logic;
	FA1854 : full_adder port map (N4_15_40,N5_0_40,N5_1_40,N6_0_40,N6_1_41);
-- In matrix 5 adding FA to column 40 
	-- signal N6_2_40 : std_logic;
	-- signal N6_3_41 : std_logic;
	FA1855 : full_adder port map (N5_2_40,N5_3_40,N5_4_40,N6_2_40,N6_3_41);
-- In matrix 5 adding FA to column 40 
	-- signal N6_4_40 : std_logic;
	-- signal N6_5_41 : std_logic;
	FA1856 : full_adder port map (N5_5_40,N5_6_40,N5_7_40,N6_4_40,N6_5_41);
-- In matrix 5 adding FA to column 41 
	-- signal N6_0_41 : std_logic;
	-- signal N6_1_42 : std_logic;
	FA1857 : full_adder port map (N4_15_41,N5_0_41,N5_1_41,N6_0_41,N6_1_42);
-- In matrix 5 adding FA to column 41 
	-- signal N6_2_41 : std_logic;
	-- signal N6_3_42 : std_logic;
	FA1858 : full_adder port map (N5_2_41,N5_3_41,N5_4_41,N6_2_41,N6_3_42);
-- In matrix 5 adding FA to column 41 
	-- signal N6_4_41 : std_logic;
	-- signal N6_5_42 : std_logic;
	FA1859 : full_adder port map (N5_5_41,N5_6_41,N5_7_41,N6_4_41,N6_5_42);
-- In matrix 5 adding FA to column 42 
	-- signal N6_0_42 : std_logic;
	-- signal N6_1_43 : std_logic;
	FA1860 : full_adder port map (N4_15_42,N5_0_42,N5_1_42,N6_0_42,N6_1_43);
-- In matrix 5 adding FA to column 42 
	-- signal N6_2_42 : std_logic;
	-- signal N6_3_43 : std_logic;
	FA1861 : full_adder port map (N5_2_42,N5_3_42,N5_4_42,N6_2_42,N6_3_43);
-- In matrix 5 adding FA to column 42 
	-- signal N6_4_42 : std_logic;
	-- signal N6_5_43 : std_logic;
	FA1862 : full_adder port map (N5_5_42,N5_6_42,N5_7_42,N6_4_42,N6_5_43);
-- In matrix 5 adding FA to column 43 
	-- signal N6_0_43 : std_logic;
	-- signal N6_1_44 : std_logic;
	FA1863 : full_adder port map (N4_15_43,N5_0_43,N5_1_43,N6_0_43,N6_1_44);
-- In matrix 5 adding FA to column 43 
	-- signal N6_2_43 : std_logic;
	-- signal N6_3_44 : std_logic;
	FA1864 : full_adder port map (N5_2_43,N5_3_43,N5_4_43,N6_2_43,N6_3_44);
-- In matrix 5 adding FA to column 43 
	-- signal N6_4_43 : std_logic;
	-- signal N6_5_44 : std_logic;
	FA1865 : full_adder port map (N5_5_43,N5_6_43,N5_7_43,N6_4_43,N6_5_44);
-- In matrix 5 adding FA to column 44 
	-- signal N6_0_44 : std_logic;
	-- signal N6_1_45 : std_logic;
	FA1866 : full_adder port map (N4_15_44,N5_0_44,N5_1_44,N6_0_44,N6_1_45);
-- In matrix 5 adding FA to column 44 
	-- signal N6_2_44 : std_logic;
	-- signal N6_3_45 : std_logic;
	FA1867 : full_adder port map (N5_2_44,N5_3_44,N5_4_44,N6_2_44,N6_3_45);
-- In matrix 5 adding FA to column 44 
	-- signal N6_4_44 : std_logic;
	-- signal N6_5_45 : std_logic;
	FA1868 : full_adder port map (N5_5_44,N5_6_44,N5_7_44,N6_4_44,N6_5_45);
-- In matrix 5 adding FA to column 45 
	-- signal N6_0_45 : std_logic;
	-- signal N6_1_46 : std_logic;
	FA1869 : full_adder port map (N4_15_45,N5_0_45,N5_1_45,N6_0_45,N6_1_46);
-- In matrix 5 adding FA to column 45 
	-- signal N6_2_45 : std_logic;
	-- signal N6_3_46 : std_logic;
	FA1870 : full_adder port map (N5_2_45,N5_3_45,N5_4_45,N6_2_45,N6_3_46);
-- In matrix 5 adding FA to column 45 
	-- signal N6_4_45 : std_logic;
	-- signal N6_5_46 : std_logic;
	FA1871 : full_adder port map (N5_5_45,N5_6_45,N5_7_45,N6_4_45,N6_5_46);
-- In matrix 5 adding FA to column 46 
	-- signal N6_0_46 : std_logic;
	-- signal N6_1_47 : std_logic;
	FA1872 : full_adder port map (N4_15_46,N5_0_46,N5_1_46,N6_0_46,N6_1_47);
-- In matrix 5 adding FA to column 46 
	-- signal N6_2_46 : std_logic;
	-- signal N6_3_47 : std_logic;
	FA1873 : full_adder port map (N5_2_46,N5_3_46,N5_4_46,N6_2_46,N6_3_47);
-- In matrix 5 adding FA to column 46 
	-- signal N6_4_46 : std_logic;
	-- signal N6_5_47 : std_logic;
	FA1874 : full_adder port map (N5_5_46,N5_6_46,N5_7_46,N6_4_46,N6_5_47);
-- In matrix 5 adding FA to column 47 
	-- signal N6_0_47 : std_logic;
	-- signal N6_1_48 : std_logic;
	FA1875 : full_adder port map (N4_15_47,N5_0_47,N5_1_47,N6_0_47,N6_1_48);
-- In matrix 5 adding FA to column 47 
	-- signal N6_2_47 : std_logic;
	-- signal N6_3_48 : std_logic;
	FA1876 : full_adder port map (N5_2_47,N5_3_47,N5_4_47,N6_2_47,N6_3_48);
-- In matrix 5 adding FA to column 47 
	-- signal N6_4_47 : std_logic;
	-- signal N6_5_48 : std_logic;
	FA1877 : full_adder port map (N5_5_47,N5_6_47,N5_7_47,N6_4_47,N6_5_48);
-- In matrix 5 adding FA to column 48 
	-- signal N6_0_48 : std_logic;
	-- signal N6_1_49 : std_logic;
	FA1878 : full_adder port map (N4_15_48,N5_0_48,N5_1_48,N6_0_48,N6_1_49);
-- In matrix 5 adding FA to column 48 
	-- signal N6_2_48 : std_logic;
	-- signal N6_3_49 : std_logic;
	FA1879 : full_adder port map (N5_2_48,N5_3_48,N5_4_48,N6_2_48,N6_3_49);
-- In matrix 5 adding FA to column 48 
	-- signal N6_4_48 : std_logic;
	-- signal N6_5_49 : std_logic;
	FA1880 : full_adder port map (N5_5_48,N5_6_48,N5_7_48,N6_4_48,N6_5_49);
-- In matrix 5 adding FA to column 49 
	-- signal N6_0_49 : std_logic;
	-- signal N6_1_50 : std_logic;
	FA1881 : full_adder port map (N4_15_49,N5_0_49,N5_1_49,N6_0_49,N6_1_50);
-- In matrix 5 adding FA to column 49 
	-- signal N6_2_49 : std_logic;
	-- signal N6_3_50 : std_logic;
	FA1882 : full_adder port map (N5_2_49,N5_3_49,N5_4_49,N6_2_49,N6_3_50);
-- In matrix 5 adding FA to column 49 
	-- signal N6_4_49 : std_logic;
	-- signal N6_5_50 : std_logic;
	FA1883 : full_adder port map (N5_5_49,N5_6_49,N5_7_49,N6_4_49,N6_5_50);
-- In matrix 5 adding FA to column 50 
	-- signal N6_0_50 : std_logic;
	-- signal N6_1_51 : std_logic;
	FA1884 : full_adder port map (N4_15_50,N5_0_50,N5_1_50,N6_0_50,N6_1_51);
-- In matrix 5 adding FA to column 50 
	-- signal N6_2_50 : std_logic;
	-- signal N6_3_51 : std_logic;
	FA1885 : full_adder port map (N5_2_50,N5_3_50,N5_4_50,N6_2_50,N6_3_51);
-- In matrix 5 adding FA to column 50 
	-- signal N6_4_50 : std_logic;
	-- signal N6_5_51 : std_logic;
	FA1886 : full_adder port map (N5_5_50,N5_6_50,N5_7_50,N6_4_50,N6_5_51);
-- In matrix 5 adding FA to column 51 
	-- signal N6_0_51 : std_logic;
	-- signal N6_1_52 : std_logic;
	FA1887 : full_adder port map (N4_15_51,N5_0_51,N5_1_51,N6_0_51,N6_1_52);
-- In matrix 5 adding FA to column 51 
	-- signal N6_2_51 : std_logic;
	-- signal N6_3_52 : std_logic;
	FA1888 : full_adder port map (N5_2_51,N5_3_51,N5_4_51,N6_2_51,N6_3_52);
-- In matrix 5 adding FA to column 51 
	-- signal N6_4_51 : std_logic;
	-- signal N6_5_52 : std_logic;
	FA1889 : full_adder port map (N5_5_51,N5_6_51,N5_7_51,N6_4_51,N6_5_52);
-- In matrix 5 adding FA to column 52 
	-- signal N6_0_52 : std_logic;
	-- signal N6_1_53 : std_logic;
	FA1890 : full_adder port map (N4_15_52,N5_0_52,N5_1_52,N6_0_52,N6_1_53);
-- In matrix 5 adding FA to column 52 
	-- signal N6_2_52 : std_logic;
	-- signal N6_3_53 : std_logic;
	FA1891 : full_adder port map (N5_2_52,N5_3_52,N5_4_52,N6_2_52,N6_3_53);
-- In matrix 5 adding FA to column 52 
	-- signal N6_4_52 : std_logic;
	-- signal N6_5_53 : std_logic;
	FA1892 : full_adder port map (N5_5_52,N5_6_52,N5_7_52,N6_4_52,N6_5_53);
-- In matrix 5 adding FA to column 53 
	-- signal N6_0_53 : std_logic;
	-- signal N6_1_54 : std_logic;
	FA1893 : full_adder port map (N4_15_53,N5_0_53,N5_1_53,N6_0_53,N6_1_54);
-- In matrix 5 adding FA to column 53 
	-- signal N6_2_53 : std_logic;
	-- signal N6_3_54 : std_logic;
	FA1894 : full_adder port map (N5_2_53,N5_3_53,N5_4_53,N6_2_53,N6_3_54);
-- In matrix 5 adding FA to column 53 
	-- signal N6_4_53 : std_logic;
	-- signal N6_5_54 : std_logic;
	FA1895 : full_adder port map (N5_5_53,N5_6_53,N5_7_53,N6_4_53,N6_5_54);
-- In matrix 5 adding FA to column 54 
	-- signal N6_0_54 : std_logic;
	-- signal N6_1_55 : std_logic;
	FA1896 : full_adder port map (N4_15_54,N5_0_54,N5_1_54,N6_0_54,N6_1_55);
-- In matrix 5 adding FA to column 54 
	-- signal N6_2_54 : std_logic;
	-- signal N6_3_55 : std_logic;
	FA1897 : full_adder port map (N5_2_54,N5_3_54,N5_4_54,N6_2_54,N6_3_55);
-- In matrix 5 adding FA to column 54 
	-- signal N6_4_54 : std_logic;
	-- signal N6_5_55 : std_logic;
	FA1898 : full_adder port map (N5_5_54,N5_6_54,N5_7_54,N6_4_54,N6_5_55);
-- In matrix 5 adding FA to column 55 
	-- signal N6_0_55 : std_logic;
	-- signal N6_1_56 : std_logic;
	FA1899 : full_adder port map (N4_15_55,N5_0_55,N5_1_55,N6_0_55,N6_1_56);
-- In matrix 5 adding FA to column 55 
	-- signal N6_2_55 : std_logic;
	-- signal N6_3_56 : std_logic;
	FA1900 : full_adder port map (N5_2_55,N5_3_55,N5_4_55,N6_2_55,N6_3_56);
-- In matrix 5 adding FA to column 55 
	-- signal N6_4_55 : std_logic;
	-- signal N6_5_56 : std_logic;
	FA1901 : full_adder port map (N5_5_55,N5_6_55,N5_7_55,N6_4_55,N6_5_56);
-- In matrix 5 adding FA to column 56 
	-- signal N6_0_56 : std_logic;
	-- signal N6_1_57 : std_logic;
	FA1902 : full_adder port map (N4_15_56,N5_0_56,N5_1_56,N6_0_56,N6_1_57);
-- In matrix 5 adding FA to column 56 
	-- signal N6_2_56 : std_logic;
	-- signal N6_3_57 : std_logic;
	FA1903 : full_adder port map (N5_2_56,N5_3_56,N5_4_56,N6_2_56,N6_3_57);
-- In matrix 5 adding FA to column 56 
	-- signal N6_4_56 : std_logic;
	-- signal N6_5_57 : std_logic;
	FA1904 : full_adder port map (N5_5_56,N5_6_56,N5_7_56,N6_4_56,N6_5_57);
-- In matrix 5 adding FA to column 57 
	-- signal N6_0_57 : std_logic;
	-- signal N6_1_58 : std_logic;
	FA1905 : full_adder port map (N4_15_57,N5_0_57,N5_1_57,N6_0_57,N6_1_58);
-- In matrix 5 adding FA to column 57 
	-- signal N6_2_57 : std_logic;
	-- signal N6_3_58 : std_logic;
	FA1906 : full_adder port map (N5_2_57,N5_3_57,N5_4_57,N6_2_57,N6_3_58);
-- In matrix 5 adding FA to column 57 
	-- signal N6_4_57 : std_logic;
	-- signal N6_5_58 : std_logic;
	FA1907 : full_adder port map (N5_5_57,N5_6_57,N5_7_57,N6_4_57,N6_5_58);
-- In matrix 5 adding FA to column 58 
	-- signal N6_0_58 : std_logic;
	-- signal N6_1_59 : std_logic;
	FA1908 : full_adder port map (N4_15_58,N5_0_58,N5_1_58,N6_0_58,N6_1_59);
-- In matrix 5 adding FA to column 58 
	-- signal N6_2_58 : std_logic;
	-- signal N6_3_59 : std_logic;
	FA1909 : full_adder port map (N5_2_58,N5_3_58,N5_4_58,N6_2_58,N6_3_59);
-- In matrix 5 adding FA to column 58 
	-- signal N6_4_58 : std_logic;
	-- signal N6_5_59 : std_logic;
	FA1910 : full_adder port map (N5_5_58,N5_6_58,N5_7_58,N6_4_58,N6_5_59);
-- In matrix 5 adding FA to column 59 
	-- signal N6_0_59 : std_logic;
	-- signal N6_1_60 : std_logic;
	FA1911 : full_adder port map (N4_15_59,N5_0_59,N5_1_59,N6_0_59,N6_1_60);
-- In matrix 5 adding FA to column 59 
	-- signal N6_2_59 : std_logic;
	-- signal N6_3_60 : std_logic;
	FA1912 : full_adder port map (N5_2_59,N5_3_59,N5_4_59,N6_2_59,N6_3_60);
-- In matrix 5 adding FA to column 59 
	-- signal N6_4_59 : std_logic;
	-- signal N6_5_60 : std_logic;
	FA1913 : full_adder port map (N5_5_59,N5_6_59,N5_7_59,N6_4_59,N6_5_60);
-- In matrix 5 adding FA to column 60 
	-- signal N6_0_60 : std_logic;
	-- signal N6_1_61 : std_logic;
	FA1914 : full_adder port map (N4_15_60,N5_0_60,N5_1_60,N6_0_60,N6_1_61);
-- In matrix 5 adding FA to column 60 
	-- signal N6_2_60 : std_logic;
	-- signal N6_3_61 : std_logic;
	FA1915 : full_adder port map (N5_2_60,N5_3_60,N5_4_60,N6_2_60,N6_3_61);
-- In matrix 5 adding FA to column 60 
	-- signal N6_4_60 : std_logic;
	-- signal N6_5_61 : std_logic;
	FA1916 : full_adder port map (N5_5_60,N5_6_60,N5_7_60,N6_4_60,N6_5_61);
-- In matrix 5 adding FA to column 61 
	-- signal N6_0_61 : std_logic;
	-- signal N6_1_62 : std_logic;
	FA1917 : full_adder port map (N4_15_61,N5_0_61,N5_1_61,N6_0_61,N6_1_62);
-- In matrix 5 adding FA to column 61 
	-- signal N6_2_61 : std_logic;
	-- signal N6_3_62 : std_logic;
	FA1918 : full_adder port map (N5_2_61,N5_3_61,N5_4_61,N6_2_61,N6_3_62);
-- In matrix 5 adding FA to column 61 
	-- signal N6_4_61 : std_logic;
	-- signal N6_5_62 : std_logic;
	FA1919 : full_adder port map (N5_5_61,N5_6_61,N5_7_61,N6_4_61,N6_5_62);
-- In matrix 5 adding FA to column 62 
	-- signal N6_0_62 : std_logic;
	-- signal N6_1_63 : std_logic;
	FA1920 : full_adder port map (N4_15_62,N5_0_62,N5_1_62,N6_0_62,N6_1_63);
-- In matrix 5 adding FA to column 62 
	-- signal N6_2_62 : std_logic;
	-- signal N6_3_63 : std_logic;
	FA1921 : full_adder port map (N5_2_62,N5_3_62,N5_4_62,N6_2_62,N6_3_63);
-- In matrix 5 adding FA to column 62 
	-- signal N6_4_62 : std_logic;
	-- signal N6_5_63 : std_logic;
	FA1922 : full_adder port map (N5_5_62,N5_6_62,N5_7_62,N6_4_62,N6_5_63);
-- In matrix 5 adding FA to column 63 
	-- signal N6_0_63 : std_logic;
	-- signal N6_1_64 : std_logic;
	FA1923 : full_adder port map (N4_15_63,N5_0_63,N5_1_63,N6_0_63,N6_1_64);
-- In matrix 5 adding FA to column 63 
	-- signal N6_2_63 : std_logic;
	-- signal N6_3_64 : std_logic;
	FA1924 : full_adder port map (N5_2_63,N5_3_63,N5_4_63,N6_2_63,N6_3_64);
-- In matrix 5 adding FA to column 63 
	-- signal N6_4_63 : std_logic;
	-- signal N6_5_64 : std_logic;
	FA1925 : full_adder port map (N5_5_63,N5_6_63,N5_7_63,N6_4_63,N6_5_64);
-- In matrix 5 adding FA to column 64 
	-- signal N6_0_64 : std_logic;
	-- signal N6_1_65 : std_logic;
	FA1926 : full_adder port map (N4_15_64,N5_0_64,N5_1_64,N6_0_64,N6_1_65);
-- In matrix 5 adding FA to column 64 
	-- signal N6_2_64 : std_logic;
	-- signal N6_3_65 : std_logic;
	FA1927 : full_adder port map (N5_2_64,N5_3_64,N5_4_64,N6_2_64,N6_3_65);
-- In matrix 5 adding FA to column 64 
	-- signal N6_4_64 : std_logic;
	-- signal N6_5_65 : std_logic;
	FA1928 : full_adder port map (N5_5_64,N5_6_64,N5_7_64,N6_4_64,N6_5_65);
-- In matrix 5 adding FA to column 65 
	-- signal N6_0_65 : std_logic;
	-- signal N6_1_66 : std_logic;
	FA1929 : full_adder port map (N4_15_65,N5_0_65,N5_1_65,N6_0_65,N6_1_66);
-- In matrix 5 adding FA to column 65 
	-- signal N6_2_65 : std_logic;
	-- signal N6_3_66 : std_logic;
	FA1930 : full_adder port map (N5_2_65,N5_3_65,N5_4_65,N6_2_65,N6_3_66);
-- In matrix 5 adding FA to column 65 
	-- signal N6_4_65 : std_logic;
	-- signal N6_5_66 : std_logic;
	FA1931 : full_adder port map (N5_5_65,N5_6_65,N5_7_65,N6_4_65,N6_5_66);
-- In matrix 5 adding FA to column 66 
	-- signal N6_0_66 : std_logic;
	-- signal N6_1_67 : std_logic;
	FA1932 : full_adder port map (N4_15_66,N5_0_66,N5_1_66,N6_0_66,N6_1_67);
-- In matrix 5 adding FA to column 66 
	-- signal N6_2_66 : std_logic;
	-- signal N6_3_67 : std_logic;
	FA1933 : full_adder port map (N5_2_66,N5_3_66,N5_4_66,N6_2_66,N6_3_67);
-- In matrix 5 adding FA to column 66 
	-- signal N6_4_66 : std_logic;
	-- signal N6_5_67 : std_logic;
	FA1934 : full_adder port map (N5_5_66,N5_6_66,N5_7_66,N6_4_66,N6_5_67);
-- In matrix 5 adding FA to column 67 
	-- signal N6_0_67 : std_logic;
	-- signal N6_1_68 : std_logic;
	FA1935 : full_adder port map (N4_15_67,N5_0_67,N5_1_67,N6_0_67,N6_1_68);
-- In matrix 5 adding FA to column 67 
	-- signal N6_2_67 : std_logic;
	-- signal N6_3_68 : std_logic;
	FA1936 : full_adder port map (N5_2_67,N5_3_67,N5_4_67,N6_2_67,N6_3_68);
-- In matrix 5 adding FA to column 67 
	-- signal N6_4_67 : std_logic;
	-- signal N6_5_68 : std_logic;
	FA1937 : full_adder port map (N5_5_67,N5_6_67,N5_7_67,N6_4_67,N6_5_68);
-- In matrix 5 adding FA to column 68 
	-- signal N6_0_68 : std_logic;
	-- signal N6_1_69 : std_logic;
	FA1938 : full_adder port map (N4_15_68,N5_0_68,N5_1_68,N6_0_68,N6_1_69);
-- In matrix 5 adding FA to column 68 
	-- signal N6_2_68 : std_logic;
	-- signal N6_3_69 : std_logic;
	FA1939 : full_adder port map (N5_2_68,N5_3_68,N5_4_68,N6_2_68,N6_3_69);
-- In matrix 5 adding FA to column 68 
	-- signal N6_4_68 : std_logic;
	-- signal N6_5_69 : std_logic;
	FA1940 : full_adder port map (N5_5_68,N5_6_68,N5_7_68,N6_4_68,N6_5_69);
-- In matrix 5 adding FA to column 69 
	-- signal N6_0_69 : std_logic;
	-- signal N6_1_70 : std_logic;
	FA1941 : full_adder port map (N4_15_69,N5_0_69,N5_1_69,N6_0_69,N6_1_70);
-- In matrix 5 adding FA to column 69 
	-- signal N6_2_69 : std_logic;
	-- signal N6_3_70 : std_logic;
	FA1942 : full_adder port map (N5_2_69,N5_3_69,N5_4_69,N6_2_69,N6_3_70);
-- In matrix 5 adding FA to column 69 
	-- signal N6_4_69 : std_logic;
	-- signal N6_5_70 : std_logic;
	FA1943 : full_adder port map (N5_5_69,N5_6_69,N5_7_69,N6_4_69,N6_5_70);
-- In matrix 5 adding FA to column 70 
	-- signal N6_0_70 : std_logic;
	-- signal N6_1_71 : std_logic;
	FA1944 : full_adder port map (N4_15_70,N5_0_70,N5_1_70,N6_0_70,N6_1_71);
-- In matrix 5 adding FA to column 70 
	-- signal N6_2_70 : std_logic;
	-- signal N6_3_71 : std_logic;
	FA1945 : full_adder port map (N5_2_70,N5_3_70,N5_4_70,N6_2_70,N6_3_71);
-- In matrix 5 adding FA to column 70 
	-- signal N6_4_70 : std_logic;
	-- signal N6_5_71 : std_logic;
	FA1946 : full_adder port map (N5_5_70,N5_6_70,N5_7_70,N6_4_70,N6_5_71);
-- In matrix 5 adding FA to column 71 
	-- signal N6_0_71 : std_logic;
	-- signal N6_1_72 : std_logic;
	FA1947 : full_adder port map (N4_15_71,N5_0_71,N5_1_71,N6_0_71,N6_1_72);
-- In matrix 5 adding FA to column 71 
	-- signal N6_2_71 : std_logic;
	-- signal N6_3_72 : std_logic;
	FA1948 : full_adder port map (N5_2_71,N5_3_71,N5_4_71,N6_2_71,N6_3_72);
-- In matrix 5 adding FA to column 71 
	-- signal N6_4_71 : std_logic;
	-- signal N6_5_72 : std_logic;
	FA1949 : full_adder port map (N5_5_71,N5_6_71,N5_7_71,N6_4_71,N6_5_72);
-- In matrix 5 adding FA to column 72 
	-- signal N6_0_72 : std_logic;
	-- signal N6_1_73 : std_logic;
	FA1950 : full_adder port map (N4_15_72,N5_0_72,N5_1_72,N6_0_72,N6_1_73);
-- In matrix 5 adding FA to column 72 
	-- signal N6_2_72 : std_logic;
	-- signal N6_3_73 : std_logic;
	FA1951 : full_adder port map (N5_2_72,N5_3_72,N5_4_72,N6_2_72,N6_3_73);
-- In matrix 5 adding FA to column 72 
	-- signal N6_4_72 : std_logic;
	-- signal N6_5_73 : std_logic;
	FA1952 : full_adder port map (N5_5_72,N5_6_72,N5_7_72,N6_4_72,N6_5_73);
-- In matrix 5 adding FA to column 73 
	-- signal N6_0_73 : std_logic;
	-- signal N6_1_74 : std_logic;
	FA1953 : full_adder port map (N4_15_73,N5_0_73,N5_1_73,N6_0_73,N6_1_74);
-- In matrix 5 adding FA to column 73 
	-- signal N6_2_73 : std_logic;
	-- signal N6_3_74 : std_logic;
	FA1954 : full_adder port map (N5_2_73,N5_3_73,N5_4_73,N6_2_73,N6_3_74);
-- In matrix 5 adding FA to column 73 
	-- signal N6_4_73 : std_logic;
	-- signal N6_5_74 : std_logic;
	FA1955 : full_adder port map (N5_5_73,N5_6_73,N5_7_73,N6_4_73,N6_5_74);
-- In matrix 5 adding FA to column 74 
	-- signal N6_0_74 : std_logic;
	-- signal N6_1_75 : std_logic;
	FA1956 : full_adder port map (N4_15_74,N5_0_74,N5_1_74,N6_0_74,N6_1_75);
-- In matrix 5 adding FA to column 74 
	-- signal N6_2_74 : std_logic;
	-- signal N6_3_75 : std_logic;
	FA1957 : full_adder port map (N5_2_74,N5_3_74,N5_4_74,N6_2_74,N6_3_75);
-- In matrix 5 adding FA to column 74 
	-- signal N6_4_74 : std_logic;
	-- signal N6_5_75 : std_logic;
	FA1958 : full_adder port map (N5_5_74,N5_6_74,N5_7_74,N6_4_74,N6_5_75);
-- In matrix 5 adding FA to column 75 
	-- signal N6_0_75 : std_logic;
	-- signal N6_1_76 : std_logic;
	FA1959 : full_adder port map (N4_15_75,N5_0_75,N5_1_75,N6_0_75,N6_1_76);
-- In matrix 5 adding FA to column 75 
	-- signal N6_2_75 : std_logic;
	-- signal N6_3_76 : std_logic;
	FA1960 : full_adder port map (N5_2_75,N5_3_75,N5_4_75,N6_2_75,N6_3_76);
-- In matrix 5 adding FA to column 75 
	-- signal N6_4_75 : std_logic;
	-- signal N6_5_76 : std_logic;
	FA1961 : full_adder port map (N5_5_75,N5_6_75,N5_7_75,N6_4_75,N6_5_76);
-- In matrix 5 adding FA to column 76 
	-- signal N6_0_76 : std_logic;
	-- signal N6_1_77 : std_logic;
	FA1962 : full_adder port map (N4_15_76,N5_0_76,N5_1_76,N6_0_76,N6_1_77);
-- In matrix 5 adding FA to column 76 
	-- signal N6_2_76 : std_logic;
	-- signal N6_3_77 : std_logic;
	FA1963 : full_adder port map (N5_2_76,N5_3_76,N5_4_76,N6_2_76,N6_3_77);
-- In matrix 5 adding FA to column 76 
	-- signal N6_4_76 : std_logic;
	-- signal N6_5_77 : std_logic;
	FA1964 : full_adder port map (N5_5_76,N5_6_76,N5_7_76,N6_4_76,N6_5_77);
-- In matrix 5 adding FA to column 77 
	-- signal N6_0_77 : std_logic;
	-- signal N6_1_78 : std_logic;
	FA1965 : full_adder port map (N4_15_77,N5_0_77,N5_1_77,N6_0_77,N6_1_78);
-- In matrix 5 adding FA to column 77 
	-- signal N6_2_77 : std_logic;
	-- signal N6_3_78 : std_logic;
	FA1966 : full_adder port map (N5_2_77,N5_3_77,N5_4_77,N6_2_77,N6_3_78);
-- In matrix 5 adding FA to column 77 
	-- signal N6_4_77 : std_logic;
	-- signal N6_5_78 : std_logic;
	FA1967 : full_adder port map (N5_5_77,N5_6_77,N5_7_77,N6_4_77,N6_5_78);
-- In matrix 5 adding FA to column 78 
	-- signal N6_0_78 : std_logic;
	-- signal N6_1_79 : std_logic;
	FA1968 : full_adder port map (N4_15_78,N5_0_78,N5_1_78,N6_0_78,N6_1_79);
-- In matrix 5 adding FA to column 78 
	-- signal N6_2_78 : std_logic;
	-- signal N6_3_79 : std_logic;
	FA1969 : full_adder port map (N5_2_78,N5_3_78,N5_4_78,N6_2_78,N6_3_79);
-- In matrix 5 adding FA to column 78 
	-- signal N6_4_78 : std_logic;
	-- signal N6_5_79 : std_logic;
	FA1970 : full_adder port map (N5_5_78,N5_6_78,N5_7_78,N6_4_78,N6_5_79);
-- In matrix 5 adding FA to column 79 
	-- signal N6_0_79 : std_logic;
	-- signal N6_1_80 : std_logic;
	FA1971 : full_adder port map (N4_15_79,N5_0_79,N5_1_79,N6_0_79,N6_1_80);
-- In matrix 5 adding FA to column 79 
	-- signal N6_2_79 : std_logic;
	-- signal N6_3_80 : std_logic;
	FA1972 : full_adder port map (N5_2_79,N5_3_79,N5_4_79,N6_2_79,N6_3_80);
-- In matrix 5 adding FA to column 79 
	-- signal N6_4_79 : std_logic;
	-- signal N6_5_80 : std_logic;
	FA1973 : full_adder port map (N5_5_79,N5_6_79,N5_7_79,N6_4_79,N6_5_80);
-- In matrix 5 adding FA to column 80 
	-- signal N6_0_80 : std_logic;
	-- signal N6_1_81 : std_logic;
	FA1974 : full_adder port map (N4_15_80,N5_0_80,N5_1_80,N6_0_80,N6_1_81);
-- In matrix 5 adding FA to column 80 
	-- signal N6_2_80 : std_logic;
	-- signal N6_3_81 : std_logic;
	FA1975 : full_adder port map (N5_2_80,N5_3_80,N5_4_80,N6_2_80,N6_3_81);
-- In matrix 5 adding FA to column 80 
	-- signal N6_4_80 : std_logic;
	-- signal N6_5_81 : std_logic;
	FA1976 : full_adder port map (N5_5_80,N5_6_80,N5_7_80,N6_4_80,N6_5_81);
-- In matrix 5 adding FA to column 81 
	-- signal N6_0_81 : std_logic;
	-- signal N6_1_82 : std_logic;
	FA1977 : full_adder port map (N4_15_81,N5_0_81,N5_1_81,N6_0_81,N6_1_82);
-- In matrix 5 adding FA to column 81 
	-- signal N6_2_81 : std_logic;
	-- signal N6_3_82 : std_logic;
	FA1978 : full_adder port map (N5_2_81,N5_3_81,N5_4_81,N6_2_81,N6_3_82);
-- In matrix 5 adding FA to column 81 
	-- signal N6_4_81 : std_logic;
	-- signal N6_5_82 : std_logic;
	FA1979 : full_adder port map (N5_5_81,N5_6_81,N5_7_81,N6_4_81,N6_5_82);
-- In matrix 5 adding FA to column 82 
	-- signal N6_0_82 : std_logic;
	-- signal N6_1_83 : std_logic;
	FA1980 : full_adder port map (N4_15_82,N5_0_82,N5_1_82,N6_0_82,N6_1_83);
-- In matrix 5 adding FA to column 82 
	-- signal N6_2_82 : std_logic;
	-- signal N6_3_83 : std_logic;
	FA1981 : full_adder port map (N5_2_82,N5_3_82,N5_4_82,N6_2_82,N6_3_83);
-- In matrix 5 adding FA to column 82 
	-- signal N6_4_82 : std_logic;
	-- signal N6_5_83 : std_logic;
	FA1982 : full_adder port map (N5_5_82,N5_6_82,N5_7_82,N6_4_82,N6_5_83);
-- In matrix 5 adding FA to column 83 
	-- signal N6_0_83 : std_logic;
	-- signal N6_1_84 : std_logic;
	FA1983 : full_adder port map (N4_15_83,N5_0_83,N5_1_83,N6_0_83,N6_1_84);
-- In matrix 5 adding FA to column 83 
	-- signal N6_2_83 : std_logic;
	-- signal N6_3_84 : std_logic;
	FA1984 : full_adder port map (N5_2_83,N5_3_83,N5_4_83,N6_2_83,N6_3_84);
-- In matrix 5 adding FA to column 83 
	-- signal N6_4_83 : std_logic;
	-- signal N6_5_84 : std_logic;
	FA1985 : full_adder port map (N5_5_83,N5_6_83,N5_7_83,N6_4_83,N6_5_84);
-- In matrix 5 adding FA to column 84 
	-- signal N6_0_84 : std_logic;
	-- signal N6_1_85 : std_logic;
	FA1986 : full_adder port map (N4_13_84,N5_0_84,N5_1_84,N6_0_84,N6_1_85);
-- In matrix 5 adding FA to column 84 
	-- signal N6_2_84 : std_logic;
	-- signal N6_3_85 : std_logic;
	FA1987 : full_adder port map (N5_2_84,N5_3_84,N5_4_84,N6_2_84,N6_3_85);
-- In matrix 5 adding FA to column 84 
	-- signal N6_4_84 : std_logic;
	-- signal N6_5_85 : std_logic;
	FA1988 : full_adder port map (N5_5_84,N5_6_84,N5_7_84,N6_4_84,N6_5_85);
-- In matrix 5 adding FA to column 85 
	-- signal N6_0_85 : std_logic;
	-- signal N6_1_86 : std_logic;
	FA1989 : full_adder port map (N4_11_85,N5_0_85,N5_1_85,N6_0_85,N6_1_86);
-- In matrix 5 adding FA to column 85 
	-- signal N6_2_85 : std_logic;
	-- signal N6_3_86 : std_logic;
	FA1990 : full_adder port map (N5_2_85,N5_3_85,N5_4_85,N6_2_85,N6_3_86);
-- In matrix 5 adding FA to column 85 
	-- signal N6_4_85 : std_logic;
	-- signal N6_5_86 : std_logic;
	FA1991 : full_adder port map (N5_5_85,N5_6_85,N5_7_85,N6_4_85,N6_5_86);
-- In matrix 5 adding FA to column 86 
	-- signal N6_0_86 : std_logic;
	-- signal N6_1_87 : std_logic;
	FA1992 : full_adder port map (N4_9_86,N5_0_86,N5_1_86,N6_0_86,N6_1_87);
-- In matrix 5 adding FA to column 86 
	-- signal N6_2_86 : std_logic;
	-- signal N6_3_87 : std_logic;
	FA1993 : full_adder port map (N5_2_86,N5_3_86,N5_4_86,N6_2_86,N6_3_87);
-- In matrix 5 adding FA to column 86 
	-- signal N6_4_86 : std_logic;
	-- signal N6_5_87 : std_logic;
	FA1994 : full_adder port map (N5_5_86,N5_6_86,N5_7_86,N6_4_86,N6_5_87);
-- In matrix 5 adding FA to column 87 
	-- signal N6_0_87 : std_logic;
	-- signal N6_1_88 : std_logic;
	FA1995 : full_adder port map (N4_7_87,N5_0_87,N5_1_87,N6_0_87,N6_1_88);
-- In matrix 5 adding FA to column 87 
	-- signal N6_2_87 : std_logic;
	-- signal N6_3_88 : std_logic;
	FA1996 : full_adder port map (N5_2_87,N5_3_87,N5_4_87,N6_2_87,N6_3_88);
-- In matrix 5 adding FA to column 87 
	-- signal N6_4_87 : std_logic;
	-- signal N6_5_88 : std_logic;
	FA1997 : full_adder port map (N5_5_87,N5_6_87,N5_7_87,N6_4_87,N6_5_88);
-- In matrix 5 adding FA to column 88 
	-- signal N6_0_88 : std_logic;
	-- signal N6_1_89 : std_logic;
	FA1998 : full_adder port map (N4_5_88,N5_0_88,N5_1_88,N6_0_88,N6_1_89);
-- In matrix 5 adding FA to column 88 
	-- signal N6_2_88 : std_logic;
	-- signal N6_3_89 : std_logic;
	FA1999 : full_adder port map (N5_2_88,N5_3_88,N5_4_88,N6_2_88,N6_3_89);
-- In matrix 5 adding FA to column 88 
	-- signal N6_4_88 : std_logic;
	-- signal N6_5_89 : std_logic;
	FA2000 : full_adder port map (N5_5_88,N5_6_88,N5_7_88,N6_4_88,N6_5_89);
-- In matrix 5 adding FA to column 89 
	-- signal N6_0_89 : std_logic;
	-- signal N6_1_90 : std_logic;
	FA2001 : full_adder port map (N4_3_89,N5_0_89,N5_1_89,N6_0_89,N6_1_90);
-- In matrix 5 adding FA to column 89 
	-- signal N6_2_89 : std_logic;
	-- signal N6_3_90 : std_logic;
	FA2002 : full_adder port map (N5_2_89,N5_3_89,N5_4_89,N6_2_89,N6_3_90);
-- In matrix 5 adding FA to column 89 
	-- signal N6_4_89 : std_logic;
	-- signal N6_5_90 : std_logic;
	FA2003 : full_adder port map (N5_5_89,N5_6_89,N5_7_89,N6_4_89,N6_5_90);
-- In matrix 5 adding FA to column 90 
	-- signal N6_0_90 : std_logic;
	-- signal N6_1_91 : std_logic;
	FA2004 : full_adder port map (N4_1_90,N5_0_90,N5_1_90,N6_0_90,N6_1_91);
-- In matrix 5 adding FA to column 90 
	-- signal N6_2_90 : std_logic;
	-- signal N6_3_91 : std_logic;
	FA2005 : full_adder port map (N5_2_90,N5_3_90,N5_4_90,N6_2_90,N6_3_91);
-- In matrix 5 adding FA to column 90 
	-- signal N6_4_90 : std_logic;
	-- signal N6_5_91 : std_logic;
	FA2006 : full_adder port map (N5_5_90,N5_6_90,N5_7_90,N6_4_90,N6_5_91);
-- In matrix 5 adding FA to column 91 
	-- signal N6_0_91 : std_logic;
	-- signal N6_1_92 : std_logic;
	FA2007 : full_adder port map (N0_51_91,N0_52_91,N5_0_91,N6_0_91,N6_1_92);
-- In matrix 5 adding FA to column 91 
	-- signal N6_2_91 : std_logic;
	-- signal N6_3_92 : std_logic;
	FA2008 : full_adder port map (N5_1_91,N5_2_91,N5_3_91,N6_2_91,N6_3_92);
-- In matrix 5 adding FA to column 91 
	-- signal N6_4_91 : std_logic;
	-- signal N6_5_92 : std_logic;
	FA2009 : full_adder port map (N5_4_91,N5_5_91,N5_6_91,N6_4_91,N6_5_92);
-- In matrix 5 adding FA to column 92 
	-- signal N6_0_92 : std_logic;
	-- signal N6_1_93 : std_logic;
	FA2010 : full_adder port map (N0_49_92,N0_50_92,N0_51_92,N6_0_92,N6_1_93);
-- In matrix 5 adding FA to column 92 
	-- signal N6_2_92 : std_logic;
	-- signal N6_3_93 : std_logic;
	FA2011 : full_adder port map (N0_52_92,N5_0_92,N5_1_92,N6_2_92,N6_3_93);
-- In matrix 5 adding FA to column 92 
	-- signal N6_4_92 : std_logic;
	-- signal N6_5_93 : std_logic;
	FA2012 : full_adder port map (N5_2_92,N5_3_92,N5_4_92,N6_4_92,N6_5_93);
-- In matrix 5 adding FA to column 93 
	-- signal N6_0_93 : std_logic;
	-- signal N6_1_94 : std_logic;
	FA2013 : full_adder port map (N0_47_93,N0_48_93,N0_49_93,N6_0_93,N6_1_94);
-- In matrix 5 adding FA to column 93 
	-- signal N6_2_93 : std_logic;
	-- signal N6_3_94 : std_logic;
	FA2014 : full_adder port map (N0_50_93,N0_51_93,N0_52_93,N6_2_93,N6_3_94);
-- In matrix 5 adding FA to column 93 
	-- signal N6_4_93 : std_logic;
	-- signal N6_5_94 : std_logic;
	FA2015 : full_adder port map (N5_0_93,N5_1_93,N5_2_93,N6_4_93,N6_5_94);
-- In matrix 5 adding FA to column 94 
	-- signal N6_0_94 : std_logic;
	-- signal N6_1_95 : std_logic;
	FA2016 : full_adder port map (N0_45_94,N0_46_94,N0_47_94,N6_0_94,N6_1_95);
-- In matrix 5 adding FA to column 94 
	-- signal N6_2_94 : std_logic;
	-- signal N6_3_95 : std_logic;
	FA2017 : full_adder port map (N0_48_94,N0_49_94,N0_50_94,N6_2_94,N6_3_95);
-- In matrix 5 adding FA to column 94 
	-- signal N6_4_94 : std_logic;
	-- signal N6_5_95 : std_logic;
	FA2018 : full_adder port map (N0_51_94,N0_52_94,N5_0_94,N6_4_94,N6_5_95);
-- In matrix 5 adding FA to column 95 
	-- signal N6_0_95 : std_logic;
	-- signal N6_1_96 : std_logic;
	FA2019 : full_adder port map (N0_43_95,N0_44_95,N0_45_95,N6_0_95,N6_1_96);
-- In matrix 5 adding FA to column 95 
	-- signal N6_2_95 : std_logic;
	-- signal N6_3_96 : std_logic;
	FA2020 : full_adder port map (N0_46_95,N0_47_95,N0_48_95,N6_2_95,N6_3_96);
-- In matrix 5 adding FA to column 95 
	-- signal N6_4_95 : std_logic;
	-- signal N6_5_96 : std_logic;
	FA2021 : full_adder port map (N0_49_95,N0_50_95,N0_51_95,N6_4_95,N6_5_96);
-- In matrix 5 adding FA to column 96 
	-- signal N6_0_96 : std_logic;
	-- signal N6_1_97 : std_logic;
	FA2022 : full_adder port map (N0_44_96,N0_45_96,N0_46_96,N6_0_96,N6_1_97);
-- In matrix 5 adding FA to column 96 
	-- signal N6_2_96 : std_logic;
	-- signal N6_3_97 : std_logic;
	FA2023 : full_adder port map (N0_47_96,N0_48_96,N0_49_96,N6_2_96,N6_3_97);
-- In matrix 5 adding FA to column 97 
	-- signal N6_0_97 : std_logic;
	-- signal N6_1_98 : std_logic;
	FA2024 : full_adder port map (N0_45_97,N0_46_97,N0_47_97,N6_0_97,N6_1_98);
	-- Elements from matrix 6 
-- In matrix 6 adding HA to column 6 
	-- signal N7_0_6 : std_logic;
	-- signal N7_1_7 : std_logic;
	HA47 : half_adder port map (N0_0_6,N0_1_6,N7_0_6,N7_1_7);
-- In matrix 6 adding FA to column 7 
	-- signal N7_0_7 : std_logic;
	-- signal N7_1_8 : std_logic;
	FA2025 : full_adder port map (N0_0_7,N0_1_7,N0_2_7,N7_0_7,N7_1_8);
-- In matrix 6 adding HA to column 7 
	-- signal N7_2_7 : std_logic;
	-- signal N7_3_8 : std_logic;
	HA48 : half_adder port map (N0_3_7,N0_4_7,N7_2_7,N7_3_8);
-- In matrix 6 adding FA to column 8 
	-- signal N7_0_8 : std_logic;
	-- signal N7_1_9 : std_logic;
	FA2026 : full_adder port map (N0_2_8,N0_3_8,N0_4_8,N7_0_8,N7_1_9);
-- In matrix 6 adding FA to column 8 
	-- signal N7_2_8 : std_logic;
	-- signal N7_3_9 : std_logic;
	FA2027 : full_adder port map (N0_5_8,N0_6_8,N0_7_8,N7_2_8,N7_3_9);
-- In matrix 6 adding FA to column 9 
	-- signal N7_0_9 : std_logic;
	-- signal N7_1_10 : std_logic;
	FA2028 : full_adder port map (N0_5_9,N0_6_9,N0_7_9,N7_0_9,N7_1_10);
-- In matrix 6 adding FA to column 9 
	-- signal N7_2_9 : std_logic;
	-- signal N7_3_10 : std_logic;
	FA2029 : full_adder port map (N0_8_9,N0_9_9,N6_0_9,N7_2_9,N7_3_10);
-- In matrix 6 adding FA to column 10 
	-- signal N7_0_10 : std_logic;
	-- signal N7_1_11 : std_logic;
	FA2030 : full_adder port map (N0_8_10,N0_9_10,N0_10_10,N7_0_10,N7_1_11);
-- In matrix 6 adding FA to column 10 
	-- signal N7_2_10 : std_logic;
	-- signal N7_3_11 : std_logic;
	FA2031 : full_adder port map (N6_0_10,N6_1_10,N6_2_10,N7_2_10,N7_3_11);
-- In matrix 6 adding FA to column 11 
	-- signal N7_0_11 : std_logic;
	-- signal N7_1_12 : std_logic;
	FA2032 : full_adder port map (N0_11_11,N5_0_11,N6_0_11,N7_0_11,N7_1_12);
-- In matrix 6 adding FA to column 11 
	-- signal N7_2_11 : std_logic;
	-- signal N7_3_12 : std_logic;
	FA2033 : full_adder port map (N6_1_11,N6_2_11,N6_3_11,N7_2_11,N7_3_12);
-- In matrix 6 adding FA to column 12 
	-- signal N7_0_12 : std_logic;
	-- signal N7_1_13 : std_logic;
	FA2034 : full_adder port map (N5_1_12,N5_2_12,N6_0_12,N7_0_12,N7_1_13);
-- In matrix 6 adding FA to column 12 
	-- signal N7_2_12 : std_logic;
	-- signal N7_3_13 : std_logic;
	FA2035 : full_adder port map (N6_1_12,N6_2_12,N6_3_12,N7_2_12,N7_3_13);
-- In matrix 6 adding FA to column 13 
	-- signal N7_0_13 : std_logic;
	-- signal N7_1_14 : std_logic;
	FA2036 : full_adder port map (N5_3_13,N5_4_13,N6_0_13,N7_0_13,N7_1_14);
-- In matrix 6 adding FA to column 13 
	-- signal N7_2_13 : std_logic;
	-- signal N7_3_14 : std_logic;
	FA2037 : full_adder port map (N6_1_13,N6_2_13,N6_3_13,N7_2_13,N7_3_14);
-- In matrix 6 adding FA to column 14 
	-- signal N7_0_14 : std_logic;
	-- signal N7_1_15 : std_logic;
	FA2038 : full_adder port map (N5_5_14,N5_6_14,N6_0_14,N7_0_14,N7_1_15);
-- In matrix 6 adding FA to column 14 
	-- signal N7_2_14 : std_logic;
	-- signal N7_3_15 : std_logic;
	FA2039 : full_adder port map (N6_1_14,N6_2_14,N6_3_14,N7_2_14,N7_3_15);
-- In matrix 6 adding FA to column 15 
	-- signal N7_0_15 : std_logic;
	-- signal N7_1_16 : std_logic;
	FA2040 : full_adder port map (N5_7_15,N5_8_15,N6_0_15,N7_0_15,N7_1_16);
-- In matrix 6 adding FA to column 15 
	-- signal N7_2_15 : std_logic;
	-- signal N7_3_16 : std_logic;
	FA2041 : full_adder port map (N6_1_15,N6_2_15,N6_3_15,N7_2_15,N7_3_16);
-- In matrix 6 adding FA to column 16 
	-- signal N7_0_16 : std_logic;
	-- signal N7_1_17 : std_logic;
	FA2042 : full_adder port map (N5_8_16,N5_9_16,N6_0_16,N7_0_16,N7_1_17);
-- In matrix 6 adding FA to column 16 
	-- signal N7_2_16 : std_logic;
	-- signal N7_3_17 : std_logic;
	FA2043 : full_adder port map (N6_1_16,N6_2_16,N6_3_16,N7_2_16,N7_3_17);
-- In matrix 6 adding FA to column 17 
	-- signal N7_0_17 : std_logic;
	-- signal N7_1_18 : std_logic;
	FA2044 : full_adder port map (N5_8_17,N5_9_17,N6_0_17,N7_0_17,N7_1_18);
-- In matrix 6 adding FA to column 17 
	-- signal N7_2_17 : std_logic;
	-- signal N7_3_18 : std_logic;
	FA2045 : full_adder port map (N6_1_17,N6_2_17,N6_3_17,N7_2_17,N7_3_18);
-- In matrix 6 adding FA to column 18 
	-- signal N7_0_18 : std_logic;
	-- signal N7_1_19 : std_logic;
	FA2046 : full_adder port map (N5_8_18,N5_9_18,N6_0_18,N7_0_18,N7_1_19);
-- In matrix 6 adding FA to column 18 
	-- signal N7_2_18 : std_logic;
	-- signal N7_3_19 : std_logic;
	FA2047 : full_adder port map (N6_1_18,N6_2_18,N6_3_18,N7_2_18,N7_3_19);
-- In matrix 6 adding FA to column 19 
	-- signal N7_0_19 : std_logic;
	-- signal N7_1_20 : std_logic;
	FA2048 : full_adder port map (N5_8_19,N5_9_19,N6_0_19,N7_0_19,N7_1_20);
-- In matrix 6 adding FA to column 19 
	-- signal N7_2_19 : std_logic;
	-- signal N7_3_20 : std_logic;
	FA2049 : full_adder port map (N6_1_19,N6_2_19,N6_3_19,N7_2_19,N7_3_20);
-- In matrix 6 adding FA to column 20 
	-- signal N7_0_20 : std_logic;
	-- signal N7_1_21 : std_logic;
	FA2050 : full_adder port map (N5_8_20,N5_9_20,N6_0_20,N7_0_20,N7_1_21);
-- In matrix 6 adding FA to column 20 
	-- signal N7_2_20 : std_logic;
	-- signal N7_3_21 : std_logic;
	FA2051 : full_adder port map (N6_1_20,N6_2_20,N6_3_20,N7_2_20,N7_3_21);
-- In matrix 6 adding FA to column 21 
	-- signal N7_0_21 : std_logic;
	-- signal N7_1_22 : std_logic;
	FA2052 : full_adder port map (N5_8_21,N5_9_21,N6_0_21,N7_0_21,N7_1_22);
-- In matrix 6 adding FA to column 21 
	-- signal N7_2_21 : std_logic;
	-- signal N7_3_22 : std_logic;
	FA2053 : full_adder port map (N6_1_21,N6_2_21,N6_3_21,N7_2_21,N7_3_22);
-- In matrix 6 adding FA to column 22 
	-- signal N7_0_22 : std_logic;
	-- signal N7_1_23 : std_logic;
	FA2054 : full_adder port map (N5_8_22,N5_9_22,N6_0_22,N7_0_22,N7_1_23);
-- In matrix 6 adding FA to column 22 
	-- signal N7_2_22 : std_logic;
	-- signal N7_3_23 : std_logic;
	FA2055 : full_adder port map (N6_1_22,N6_2_22,N6_3_22,N7_2_22,N7_3_23);
-- In matrix 6 adding FA to column 23 
	-- signal N7_0_23 : std_logic;
	-- signal N7_1_24 : std_logic;
	FA2056 : full_adder port map (N5_8_23,N5_9_23,N6_0_23,N7_0_23,N7_1_24);
-- In matrix 6 adding FA to column 23 
	-- signal N7_2_23 : std_logic;
	-- signal N7_3_24 : std_logic;
	FA2057 : full_adder port map (N6_1_23,N6_2_23,N6_3_23,N7_2_23,N7_3_24);
-- In matrix 6 adding FA to column 24 
	-- signal N7_0_24 : std_logic;
	-- signal N7_1_25 : std_logic;
	FA2058 : full_adder port map (N5_8_24,N5_9_24,N6_0_24,N7_0_24,N7_1_25);
-- In matrix 6 adding FA to column 24 
	-- signal N7_2_24 : std_logic;
	-- signal N7_3_25 : std_logic;
	FA2059 : full_adder port map (N6_1_24,N6_2_24,N6_3_24,N7_2_24,N7_3_25);
-- In matrix 6 adding FA to column 25 
	-- signal N7_0_25 : std_logic;
	-- signal N7_1_26 : std_logic;
	FA2060 : full_adder port map (N5_8_25,N5_9_25,N6_0_25,N7_0_25,N7_1_26);
-- In matrix 6 adding FA to column 25 
	-- signal N7_2_25 : std_logic;
	-- signal N7_3_26 : std_logic;
	FA2061 : full_adder port map (N6_1_25,N6_2_25,N6_3_25,N7_2_25,N7_3_26);
-- In matrix 6 adding FA to column 26 
	-- signal N7_0_26 : std_logic;
	-- signal N7_1_27 : std_logic;
	FA2062 : full_adder port map (N5_8_26,N5_9_26,N6_0_26,N7_0_26,N7_1_27);
-- In matrix 6 adding FA to column 26 
	-- signal N7_2_26 : std_logic;
	-- signal N7_3_27 : std_logic;
	FA2063 : full_adder port map (N6_1_26,N6_2_26,N6_3_26,N7_2_26,N7_3_27);
-- In matrix 6 adding FA to column 27 
	-- signal N7_0_27 : std_logic;
	-- signal N7_1_28 : std_logic;
	FA2064 : full_adder port map (N5_8_27,N5_9_27,N6_0_27,N7_0_27,N7_1_28);
-- In matrix 6 adding FA to column 27 
	-- signal N7_2_27 : std_logic;
	-- signal N7_3_28 : std_logic;
	FA2065 : full_adder port map (N6_1_27,N6_2_27,N6_3_27,N7_2_27,N7_3_28);
-- In matrix 6 adding FA to column 28 
	-- signal N7_0_28 : std_logic;
	-- signal N7_1_29 : std_logic;
	FA2066 : full_adder port map (N5_8_28,N5_9_28,N6_0_28,N7_0_28,N7_1_29);
-- In matrix 6 adding FA to column 28 
	-- signal N7_2_28 : std_logic;
	-- signal N7_3_29 : std_logic;
	FA2067 : full_adder port map (N6_1_28,N6_2_28,N6_3_28,N7_2_28,N7_3_29);
-- In matrix 6 adding FA to column 29 
	-- signal N7_0_29 : std_logic;
	-- signal N7_1_30 : std_logic;
	FA2068 : full_adder port map (N5_8_29,N5_9_29,N6_0_29,N7_0_29,N7_1_30);
-- In matrix 6 adding FA to column 29 
	-- signal N7_2_29 : std_logic;
	-- signal N7_3_30 : std_logic;
	FA2069 : full_adder port map (N6_1_29,N6_2_29,N6_3_29,N7_2_29,N7_3_30);
-- In matrix 6 adding FA to column 30 
	-- signal N7_0_30 : std_logic;
	-- signal N7_1_31 : std_logic;
	FA2070 : full_adder port map (N5_8_30,N5_9_30,N6_0_30,N7_0_30,N7_1_31);
-- In matrix 6 adding FA to column 30 
	-- signal N7_2_30 : std_logic;
	-- signal N7_3_31 : std_logic;
	FA2071 : full_adder port map (N6_1_30,N6_2_30,N6_3_30,N7_2_30,N7_3_31);
-- In matrix 6 adding FA to column 31 
	-- signal N7_0_31 : std_logic;
	-- signal N7_1_32 : std_logic;
	FA2072 : full_adder port map (N5_8_31,N5_9_31,N6_0_31,N7_0_31,N7_1_32);
-- In matrix 6 adding FA to column 31 
	-- signal N7_2_31 : std_logic;
	-- signal N7_3_32 : std_logic;
	FA2073 : full_adder port map (N6_1_31,N6_2_31,N6_3_31,N7_2_31,N7_3_32);
-- In matrix 6 adding FA to column 32 
	-- signal N7_0_32 : std_logic;
	-- signal N7_1_33 : std_logic;
	FA2074 : full_adder port map (N5_8_32,N5_9_32,N6_0_32,N7_0_32,N7_1_33);
-- In matrix 6 adding FA to column 32 
	-- signal N7_2_32 : std_logic;
	-- signal N7_3_33 : std_logic;
	FA2075 : full_adder port map (N6_1_32,N6_2_32,N6_3_32,N7_2_32,N7_3_33);
-- In matrix 6 adding FA to column 33 
	-- signal N7_0_33 : std_logic;
	-- signal N7_1_34 : std_logic;
	FA2076 : full_adder port map (N5_8_33,N5_9_33,N6_0_33,N7_0_33,N7_1_34);
-- In matrix 6 adding FA to column 33 
	-- signal N7_2_33 : std_logic;
	-- signal N7_3_34 : std_logic;
	FA2077 : full_adder port map (N6_1_33,N6_2_33,N6_3_33,N7_2_33,N7_3_34);
-- In matrix 6 adding FA to column 34 
	-- signal N7_0_34 : std_logic;
	-- signal N7_1_35 : std_logic;
	FA2078 : full_adder port map (N5_8_34,N5_9_34,N6_0_34,N7_0_34,N7_1_35);
-- In matrix 6 adding FA to column 34 
	-- signal N7_2_34 : std_logic;
	-- signal N7_3_35 : std_logic;
	FA2079 : full_adder port map (N6_1_34,N6_2_34,N6_3_34,N7_2_34,N7_3_35);
-- In matrix 6 adding FA to column 35 
	-- signal N7_0_35 : std_logic;
	-- signal N7_1_36 : std_logic;
	FA2080 : full_adder port map (N5_8_35,N5_9_35,N6_0_35,N7_0_35,N7_1_36);
-- In matrix 6 adding FA to column 35 
	-- signal N7_2_35 : std_logic;
	-- signal N7_3_36 : std_logic;
	FA2081 : full_adder port map (N6_1_35,N6_2_35,N6_3_35,N7_2_35,N7_3_36);
-- In matrix 6 adding FA to column 36 
	-- signal N7_0_36 : std_logic;
	-- signal N7_1_37 : std_logic;
	FA2082 : full_adder port map (N5_8_36,N5_9_36,N6_0_36,N7_0_36,N7_1_37);
-- In matrix 6 adding FA to column 36 
	-- signal N7_2_36 : std_logic;
	-- signal N7_3_37 : std_logic;
	FA2083 : full_adder port map (N6_1_36,N6_2_36,N6_3_36,N7_2_36,N7_3_37);
-- In matrix 6 adding FA to column 37 
	-- signal N7_0_37 : std_logic;
	-- signal N7_1_38 : std_logic;
	FA2084 : full_adder port map (N5_8_37,N5_9_37,N6_0_37,N7_0_37,N7_1_38);
-- In matrix 6 adding FA to column 37 
	-- signal N7_2_37 : std_logic;
	-- signal N7_3_38 : std_logic;
	FA2085 : full_adder port map (N6_1_37,N6_2_37,N6_3_37,N7_2_37,N7_3_38);
-- In matrix 6 adding FA to column 38 
	-- signal N7_0_38 : std_logic;
	-- signal N7_1_39 : std_logic;
	FA2086 : full_adder port map (N5_8_38,N5_9_38,N6_0_38,N7_0_38,N7_1_39);
-- In matrix 6 adding FA to column 38 
	-- signal N7_2_38 : std_logic;
	-- signal N7_3_39 : std_logic;
	FA2087 : full_adder port map (N6_1_38,N6_2_38,N6_3_38,N7_2_38,N7_3_39);
-- In matrix 6 adding FA to column 39 
	-- signal N7_0_39 : std_logic;
	-- signal N7_1_40 : std_logic;
	FA2088 : full_adder port map (N5_8_39,N5_9_39,N6_0_39,N7_0_39,N7_1_40);
-- In matrix 6 adding FA to column 39 
	-- signal N7_2_39 : std_logic;
	-- signal N7_3_40 : std_logic;
	FA2089 : full_adder port map (N6_1_39,N6_2_39,N6_3_39,N7_2_39,N7_3_40);
-- In matrix 6 adding FA to column 40 
	-- signal N7_0_40 : std_logic;
	-- signal N7_1_41 : std_logic;
	FA2090 : full_adder port map (N5_8_40,N5_9_40,N6_0_40,N7_0_40,N7_1_41);
-- In matrix 6 adding FA to column 40 
	-- signal N7_2_40 : std_logic;
	-- signal N7_3_41 : std_logic;
	FA2091 : full_adder port map (N6_1_40,N6_2_40,N6_3_40,N7_2_40,N7_3_41);
-- In matrix 6 adding FA to column 41 
	-- signal N7_0_41 : std_logic;
	-- signal N7_1_42 : std_logic;
	FA2092 : full_adder port map (N5_8_41,N5_9_41,N6_0_41,N7_0_41,N7_1_42);
-- In matrix 6 adding FA to column 41 
	-- signal N7_2_41 : std_logic;
	-- signal N7_3_42 : std_logic;
	FA2093 : full_adder port map (N6_1_41,N6_2_41,N6_3_41,N7_2_41,N7_3_42);
-- In matrix 6 adding FA to column 42 
	-- signal N7_0_42 : std_logic;
	-- signal N7_1_43 : std_logic;
	FA2094 : full_adder port map (N5_8_42,N5_9_42,N6_0_42,N7_0_42,N7_1_43);
-- In matrix 6 adding FA to column 42 
	-- signal N7_2_42 : std_logic;
	-- signal N7_3_43 : std_logic;
	FA2095 : full_adder port map (N6_1_42,N6_2_42,N6_3_42,N7_2_42,N7_3_43);
-- In matrix 6 adding FA to column 43 
	-- signal N7_0_43 : std_logic;
	-- signal N7_1_44 : std_logic;
	FA2096 : full_adder port map (N5_8_43,N5_9_43,N6_0_43,N7_0_43,N7_1_44);
-- In matrix 6 adding FA to column 43 
	-- signal N7_2_43 : std_logic;
	-- signal N7_3_44 : std_logic;
	FA2097 : full_adder port map (N6_1_43,N6_2_43,N6_3_43,N7_2_43,N7_3_44);
-- In matrix 6 adding FA to column 44 
	-- signal N7_0_44 : std_logic;
	-- signal N7_1_45 : std_logic;
	FA2098 : full_adder port map (N5_8_44,N5_9_44,N6_0_44,N7_0_44,N7_1_45);
-- In matrix 6 adding FA to column 44 
	-- signal N7_2_44 : std_logic;
	-- signal N7_3_45 : std_logic;
	FA2099 : full_adder port map (N6_1_44,N6_2_44,N6_3_44,N7_2_44,N7_3_45);
-- In matrix 6 adding FA to column 45 
	-- signal N7_0_45 : std_logic;
	-- signal N7_1_46 : std_logic;
	FA2100 : full_adder port map (N5_8_45,N5_9_45,N6_0_45,N7_0_45,N7_1_46);
-- In matrix 6 adding FA to column 45 
	-- signal N7_2_45 : std_logic;
	-- signal N7_3_46 : std_logic;
	FA2101 : full_adder port map (N6_1_45,N6_2_45,N6_3_45,N7_2_45,N7_3_46);
-- In matrix 6 adding FA to column 46 
	-- signal N7_0_46 : std_logic;
	-- signal N7_1_47 : std_logic;
	FA2102 : full_adder port map (N5_8_46,N5_9_46,N6_0_46,N7_0_46,N7_1_47);
-- In matrix 6 adding FA to column 46 
	-- signal N7_2_46 : std_logic;
	-- signal N7_3_47 : std_logic;
	FA2103 : full_adder port map (N6_1_46,N6_2_46,N6_3_46,N7_2_46,N7_3_47);
-- In matrix 6 adding FA to column 47 
	-- signal N7_0_47 : std_logic;
	-- signal N7_1_48 : std_logic;
	FA2104 : full_adder port map (N5_8_47,N5_9_47,N6_0_47,N7_0_47,N7_1_48);
-- In matrix 6 adding FA to column 47 
	-- signal N7_2_47 : std_logic;
	-- signal N7_3_48 : std_logic;
	FA2105 : full_adder port map (N6_1_47,N6_2_47,N6_3_47,N7_2_47,N7_3_48);
-- In matrix 6 adding FA to column 48 
	-- signal N7_0_48 : std_logic;
	-- signal N7_1_49 : std_logic;
	FA2106 : full_adder port map (N5_8_48,N5_9_48,N6_0_48,N7_0_48,N7_1_49);
-- In matrix 6 adding FA to column 48 
	-- signal N7_2_48 : std_logic;
	-- signal N7_3_49 : std_logic;
	FA2107 : full_adder port map (N6_1_48,N6_2_48,N6_3_48,N7_2_48,N7_3_49);
-- In matrix 6 adding FA to column 49 
	-- signal N7_0_49 : std_logic;
	-- signal N7_1_50 : std_logic;
	FA2108 : full_adder port map (N5_8_49,N5_9_49,N6_0_49,N7_0_49,N7_1_50);
-- In matrix 6 adding FA to column 49 
	-- signal N7_2_49 : std_logic;
	-- signal N7_3_50 : std_logic;
	FA2109 : full_adder port map (N6_1_49,N6_2_49,N6_3_49,N7_2_49,N7_3_50);
-- In matrix 6 adding FA to column 50 
	-- signal N7_0_50 : std_logic;
	-- signal N7_1_51 : std_logic;
	FA2110 : full_adder port map (N5_8_50,N5_9_50,N6_0_50,N7_0_50,N7_1_51);
-- In matrix 6 adding FA to column 50 
	-- signal N7_2_50 : std_logic;
	-- signal N7_3_51 : std_logic;
	FA2111 : full_adder port map (N6_1_50,N6_2_50,N6_3_50,N7_2_50,N7_3_51);
-- In matrix 6 adding FA to column 51 
	-- signal N7_0_51 : std_logic;
	-- signal N7_1_52 : std_logic;
	FA2112 : full_adder port map (N5_8_51,N5_9_51,N6_0_51,N7_0_51,N7_1_52);
-- In matrix 6 adding FA to column 51 
	-- signal N7_2_51 : std_logic;
	-- signal N7_3_52 : std_logic;
	FA2113 : full_adder port map (N6_1_51,N6_2_51,N6_3_51,N7_2_51,N7_3_52);
-- In matrix 6 adding FA to column 52 
	-- signal N7_0_52 : std_logic;
	-- signal N7_1_53 : std_logic;
	FA2114 : full_adder port map (N5_8_52,N5_9_52,N6_0_52,N7_0_52,N7_1_53);
-- In matrix 6 adding FA to column 52 
	-- signal N7_2_52 : std_logic;
	-- signal N7_3_53 : std_logic;
	FA2115 : full_adder port map (N6_1_52,N6_2_52,N6_3_52,N7_2_52,N7_3_53);
-- In matrix 6 adding FA to column 53 
	-- signal N7_0_53 : std_logic;
	-- signal N7_1_54 : std_logic;
	FA2116 : full_adder port map (N5_8_53,N5_9_53,N6_0_53,N7_0_53,N7_1_54);
-- In matrix 6 adding FA to column 53 
	-- signal N7_2_53 : std_logic;
	-- signal N7_3_54 : std_logic;
	FA2117 : full_adder port map (N6_1_53,N6_2_53,N6_3_53,N7_2_53,N7_3_54);
-- In matrix 6 adding FA to column 54 
	-- signal N7_0_54 : std_logic;
	-- signal N7_1_55 : std_logic;
	FA2118 : full_adder port map (N5_8_54,N5_9_54,N6_0_54,N7_0_54,N7_1_55);
-- In matrix 6 adding FA to column 54 
	-- signal N7_2_54 : std_logic;
	-- signal N7_3_55 : std_logic;
	FA2119 : full_adder port map (N6_1_54,N6_2_54,N6_3_54,N7_2_54,N7_3_55);
-- In matrix 6 adding FA to column 55 
	-- signal N7_0_55 : std_logic;
	-- signal N7_1_56 : std_logic;
	FA2120 : full_adder port map (N5_8_55,N5_9_55,N6_0_55,N7_0_55,N7_1_56);
-- In matrix 6 adding FA to column 55 
	-- signal N7_2_55 : std_logic;
	-- signal N7_3_56 : std_logic;
	FA2121 : full_adder port map (N6_1_55,N6_2_55,N6_3_55,N7_2_55,N7_3_56);
-- In matrix 6 adding FA to column 56 
	-- signal N7_0_56 : std_logic;
	-- signal N7_1_57 : std_logic;
	FA2122 : full_adder port map (N5_8_56,N5_9_56,N6_0_56,N7_0_56,N7_1_57);
-- In matrix 6 adding FA to column 56 
	-- signal N7_2_56 : std_logic;
	-- signal N7_3_57 : std_logic;
	FA2123 : full_adder port map (N6_1_56,N6_2_56,N6_3_56,N7_2_56,N7_3_57);
-- In matrix 6 adding FA to column 57 
	-- signal N7_0_57 : std_logic;
	-- signal N7_1_58 : std_logic;
	FA2124 : full_adder port map (N5_8_57,N5_9_57,N6_0_57,N7_0_57,N7_1_58);
-- In matrix 6 adding FA to column 57 
	-- signal N7_2_57 : std_logic;
	-- signal N7_3_58 : std_logic;
	FA2125 : full_adder port map (N6_1_57,N6_2_57,N6_3_57,N7_2_57,N7_3_58);
-- In matrix 6 adding FA to column 58 
	-- signal N7_0_58 : std_logic;
	-- signal N7_1_59 : std_logic;
	FA2126 : full_adder port map (N5_8_58,N5_9_58,N6_0_58,N7_0_58,N7_1_59);
-- In matrix 6 adding FA to column 58 
	-- signal N7_2_58 : std_logic;
	-- signal N7_3_59 : std_logic;
	FA2127 : full_adder port map (N6_1_58,N6_2_58,N6_3_58,N7_2_58,N7_3_59);
-- In matrix 6 adding FA to column 59 
	-- signal N7_0_59 : std_logic;
	-- signal N7_1_60 : std_logic;
	FA2128 : full_adder port map (N5_8_59,N5_9_59,N6_0_59,N7_0_59,N7_1_60);
-- In matrix 6 adding FA to column 59 
	-- signal N7_2_59 : std_logic;
	-- signal N7_3_60 : std_logic;
	FA2129 : full_adder port map (N6_1_59,N6_2_59,N6_3_59,N7_2_59,N7_3_60);
-- In matrix 6 adding FA to column 60 
	-- signal N7_0_60 : std_logic;
	-- signal N7_1_61 : std_logic;
	FA2130 : full_adder port map (N5_8_60,N5_9_60,N6_0_60,N7_0_60,N7_1_61);
-- In matrix 6 adding FA to column 60 
	-- signal N7_2_60 : std_logic;
	-- signal N7_3_61 : std_logic;
	FA2131 : full_adder port map (N6_1_60,N6_2_60,N6_3_60,N7_2_60,N7_3_61);
-- In matrix 6 adding FA to column 61 
	-- signal N7_0_61 : std_logic;
	-- signal N7_1_62 : std_logic;
	FA2132 : full_adder port map (N5_8_61,N5_9_61,N6_0_61,N7_0_61,N7_1_62);
-- In matrix 6 adding FA to column 61 
	-- signal N7_2_61 : std_logic;
	-- signal N7_3_62 : std_logic;
	FA2133 : full_adder port map (N6_1_61,N6_2_61,N6_3_61,N7_2_61,N7_3_62);
-- In matrix 6 adding FA to column 62 
	-- signal N7_0_62 : std_logic;
	-- signal N7_1_63 : std_logic;
	FA2134 : full_adder port map (N5_8_62,N5_9_62,N6_0_62,N7_0_62,N7_1_63);
-- In matrix 6 adding FA to column 62 
	-- signal N7_2_62 : std_logic;
	-- signal N7_3_63 : std_logic;
	FA2135 : full_adder port map (N6_1_62,N6_2_62,N6_3_62,N7_2_62,N7_3_63);
-- In matrix 6 adding FA to column 63 
	-- signal N7_0_63 : std_logic;
	-- signal N7_1_64 : std_logic;
	FA2136 : full_adder port map (N5_8_63,N5_9_63,N6_0_63,N7_0_63,N7_1_64);
-- In matrix 6 adding FA to column 63 
	-- signal N7_2_63 : std_logic;
	-- signal N7_3_64 : std_logic;
	FA2137 : full_adder port map (N6_1_63,N6_2_63,N6_3_63,N7_2_63,N7_3_64);
-- In matrix 6 adding FA to column 64 
	-- signal N7_0_64 : std_logic;
	-- signal N7_1_65 : std_logic;
	FA2138 : full_adder port map (N5_8_64,N5_9_64,N6_0_64,N7_0_64,N7_1_65);
-- In matrix 6 adding FA to column 64 
	-- signal N7_2_64 : std_logic;
	-- signal N7_3_65 : std_logic;
	FA2139 : full_adder port map (N6_1_64,N6_2_64,N6_3_64,N7_2_64,N7_3_65);
-- In matrix 6 adding FA to column 65 
	-- signal N7_0_65 : std_logic;
	-- signal N7_1_66 : std_logic;
	FA2140 : full_adder port map (N5_8_65,N5_9_65,N6_0_65,N7_0_65,N7_1_66);
-- In matrix 6 adding FA to column 65 
	-- signal N7_2_65 : std_logic;
	-- signal N7_3_66 : std_logic;
	FA2141 : full_adder port map (N6_1_65,N6_2_65,N6_3_65,N7_2_65,N7_3_66);
-- In matrix 6 adding FA to column 66 
	-- signal N7_0_66 : std_logic;
	-- signal N7_1_67 : std_logic;
	FA2142 : full_adder port map (N5_8_66,N5_9_66,N6_0_66,N7_0_66,N7_1_67);
-- In matrix 6 adding FA to column 66 
	-- signal N7_2_66 : std_logic;
	-- signal N7_3_67 : std_logic;
	FA2143 : full_adder port map (N6_1_66,N6_2_66,N6_3_66,N7_2_66,N7_3_67);
-- In matrix 6 adding FA to column 67 
	-- signal N7_0_67 : std_logic;
	-- signal N7_1_68 : std_logic;
	FA2144 : full_adder port map (N5_8_67,N5_9_67,N6_0_67,N7_0_67,N7_1_68);
-- In matrix 6 adding FA to column 67 
	-- signal N7_2_67 : std_logic;
	-- signal N7_3_68 : std_logic;
	FA2145 : full_adder port map (N6_1_67,N6_2_67,N6_3_67,N7_2_67,N7_3_68);
-- In matrix 6 adding FA to column 68 
	-- signal N7_0_68 : std_logic;
	-- signal N7_1_69 : std_logic;
	FA2146 : full_adder port map (N5_8_68,N5_9_68,N6_0_68,N7_0_68,N7_1_69);
-- In matrix 6 adding FA to column 68 
	-- signal N7_2_68 : std_logic;
	-- signal N7_3_69 : std_logic;
	FA2147 : full_adder port map (N6_1_68,N6_2_68,N6_3_68,N7_2_68,N7_3_69);
-- In matrix 6 adding FA to column 69 
	-- signal N7_0_69 : std_logic;
	-- signal N7_1_70 : std_logic;
	FA2148 : full_adder port map (N5_8_69,N5_9_69,N6_0_69,N7_0_69,N7_1_70);
-- In matrix 6 adding FA to column 69 
	-- signal N7_2_69 : std_logic;
	-- signal N7_3_70 : std_logic;
	FA2149 : full_adder port map (N6_1_69,N6_2_69,N6_3_69,N7_2_69,N7_3_70);
-- In matrix 6 adding FA to column 70 
	-- signal N7_0_70 : std_logic;
	-- signal N7_1_71 : std_logic;
	FA2150 : full_adder port map (N5_8_70,N5_9_70,N6_0_70,N7_0_70,N7_1_71);
-- In matrix 6 adding FA to column 70 
	-- signal N7_2_70 : std_logic;
	-- signal N7_3_71 : std_logic;
	FA2151 : full_adder port map (N6_1_70,N6_2_70,N6_3_70,N7_2_70,N7_3_71);
-- In matrix 6 adding FA to column 71 
	-- signal N7_0_71 : std_logic;
	-- signal N7_1_72 : std_logic;
	FA2152 : full_adder port map (N5_8_71,N5_9_71,N6_0_71,N7_0_71,N7_1_72);
-- In matrix 6 adding FA to column 71 
	-- signal N7_2_71 : std_logic;
	-- signal N7_3_72 : std_logic;
	FA2153 : full_adder port map (N6_1_71,N6_2_71,N6_3_71,N7_2_71,N7_3_72);
-- In matrix 6 adding FA to column 72 
	-- signal N7_0_72 : std_logic;
	-- signal N7_1_73 : std_logic;
	FA2154 : full_adder port map (N5_8_72,N5_9_72,N6_0_72,N7_0_72,N7_1_73);
-- In matrix 6 adding FA to column 72 
	-- signal N7_2_72 : std_logic;
	-- signal N7_3_73 : std_logic;
	FA2155 : full_adder port map (N6_1_72,N6_2_72,N6_3_72,N7_2_72,N7_3_73);
-- In matrix 6 adding FA to column 73 
	-- signal N7_0_73 : std_logic;
	-- signal N7_1_74 : std_logic;
	FA2156 : full_adder port map (N5_8_73,N5_9_73,N6_0_73,N7_0_73,N7_1_74);
-- In matrix 6 adding FA to column 73 
	-- signal N7_2_73 : std_logic;
	-- signal N7_3_74 : std_logic;
	FA2157 : full_adder port map (N6_1_73,N6_2_73,N6_3_73,N7_2_73,N7_3_74);
-- In matrix 6 adding FA to column 74 
	-- signal N7_0_74 : std_logic;
	-- signal N7_1_75 : std_logic;
	FA2158 : full_adder port map (N5_8_74,N5_9_74,N6_0_74,N7_0_74,N7_1_75);
-- In matrix 6 adding FA to column 74 
	-- signal N7_2_74 : std_logic;
	-- signal N7_3_75 : std_logic;
	FA2159 : full_adder port map (N6_1_74,N6_2_74,N6_3_74,N7_2_74,N7_3_75);
-- In matrix 6 adding FA to column 75 
	-- signal N7_0_75 : std_logic;
	-- signal N7_1_76 : std_logic;
	FA2160 : full_adder port map (N5_8_75,N5_9_75,N6_0_75,N7_0_75,N7_1_76);
-- In matrix 6 adding FA to column 75 
	-- signal N7_2_75 : std_logic;
	-- signal N7_3_76 : std_logic;
	FA2161 : full_adder port map (N6_1_75,N6_2_75,N6_3_75,N7_2_75,N7_3_76);
-- In matrix 6 adding FA to column 76 
	-- signal N7_0_76 : std_logic;
	-- signal N7_1_77 : std_logic;
	FA2162 : full_adder port map (N5_8_76,N5_9_76,N6_0_76,N7_0_76,N7_1_77);
-- In matrix 6 adding FA to column 76 
	-- signal N7_2_76 : std_logic;
	-- signal N7_3_77 : std_logic;
	FA2163 : full_adder port map (N6_1_76,N6_2_76,N6_3_76,N7_2_76,N7_3_77);
-- In matrix 6 adding FA to column 77 
	-- signal N7_0_77 : std_logic;
	-- signal N7_1_78 : std_logic;
	FA2164 : full_adder port map (N5_8_77,N5_9_77,N6_0_77,N7_0_77,N7_1_78);
-- In matrix 6 adding FA to column 77 
	-- signal N7_2_77 : std_logic;
	-- signal N7_3_78 : std_logic;
	FA2165 : full_adder port map (N6_1_77,N6_2_77,N6_3_77,N7_2_77,N7_3_78);
-- In matrix 6 adding FA to column 78 
	-- signal N7_0_78 : std_logic;
	-- signal N7_1_79 : std_logic;
	FA2166 : full_adder port map (N5_8_78,N5_9_78,N6_0_78,N7_0_78,N7_1_79);
-- In matrix 6 adding FA to column 78 
	-- signal N7_2_78 : std_logic;
	-- signal N7_3_79 : std_logic;
	FA2167 : full_adder port map (N6_1_78,N6_2_78,N6_3_78,N7_2_78,N7_3_79);
-- In matrix 6 adding FA to column 79 
	-- signal N7_0_79 : std_logic;
	-- signal N7_1_80 : std_logic;
	FA2168 : full_adder port map (N5_8_79,N5_9_79,N6_0_79,N7_0_79,N7_1_80);
-- In matrix 6 adding FA to column 79 
	-- signal N7_2_79 : std_logic;
	-- signal N7_3_80 : std_logic;
	FA2169 : full_adder port map (N6_1_79,N6_2_79,N6_3_79,N7_2_79,N7_3_80);
-- In matrix 6 adding FA to column 80 
	-- signal N7_0_80 : std_logic;
	-- signal N7_1_81 : std_logic;
	FA2170 : full_adder port map (N5_8_80,N5_9_80,N6_0_80,N7_0_80,N7_1_81);
-- In matrix 6 adding FA to column 80 
	-- signal N7_2_80 : std_logic;
	-- signal N7_3_81 : std_logic;
	FA2171 : full_adder port map (N6_1_80,N6_2_80,N6_3_80,N7_2_80,N7_3_81);
-- In matrix 6 adding FA to column 81 
	-- signal N7_0_81 : std_logic;
	-- signal N7_1_82 : std_logic;
	FA2172 : full_adder port map (N5_8_81,N5_9_81,N6_0_81,N7_0_81,N7_1_82);
-- In matrix 6 adding FA to column 81 
	-- signal N7_2_81 : std_logic;
	-- signal N7_3_82 : std_logic;
	FA2173 : full_adder port map (N6_1_81,N6_2_81,N6_3_81,N7_2_81,N7_3_82);
-- In matrix 6 adding FA to column 82 
	-- signal N7_0_82 : std_logic;
	-- signal N7_1_83 : std_logic;
	FA2174 : full_adder port map (N5_8_82,N5_9_82,N6_0_82,N7_0_82,N7_1_83);
-- In matrix 6 adding FA to column 82 
	-- signal N7_2_82 : std_logic;
	-- signal N7_3_83 : std_logic;
	FA2175 : full_adder port map (N6_1_82,N6_2_82,N6_3_82,N7_2_82,N7_3_83);
-- In matrix 6 adding FA to column 83 
	-- signal N7_0_83 : std_logic;
	-- signal N7_1_84 : std_logic;
	FA2176 : full_adder port map (N5_8_83,N5_9_83,N6_0_83,N7_0_83,N7_1_84);
-- In matrix 6 adding FA to column 83 
	-- signal N7_2_83 : std_logic;
	-- signal N7_3_84 : std_logic;
	FA2177 : full_adder port map (N6_1_83,N6_2_83,N6_3_83,N7_2_83,N7_3_84);
-- In matrix 6 adding FA to column 84 
	-- signal N7_0_84 : std_logic;
	-- signal N7_1_85 : std_logic;
	FA2178 : full_adder port map (N5_8_84,N5_9_84,N6_0_84,N7_0_84,N7_1_85);
-- In matrix 6 adding FA to column 84 
	-- signal N7_2_84 : std_logic;
	-- signal N7_3_85 : std_logic;
	FA2179 : full_adder port map (N6_1_84,N6_2_84,N6_3_84,N7_2_84,N7_3_85);
-- In matrix 6 adding FA to column 85 
	-- signal N7_0_85 : std_logic;
	-- signal N7_1_86 : std_logic;
	FA2180 : full_adder port map (N5_8_85,N5_9_85,N6_0_85,N7_0_85,N7_1_86);
-- In matrix 6 adding FA to column 85 
	-- signal N7_2_85 : std_logic;
	-- signal N7_3_86 : std_logic;
	FA2181 : full_adder port map (N6_1_85,N6_2_85,N6_3_85,N7_2_85,N7_3_86);
-- In matrix 6 adding FA to column 86 
	-- signal N7_0_86 : std_logic;
	-- signal N7_1_87 : std_logic;
	FA2182 : full_adder port map (N5_8_86,N5_9_86,N6_0_86,N7_0_86,N7_1_87);
-- In matrix 6 adding FA to column 86 
	-- signal N7_2_86 : std_logic;
	-- signal N7_3_87 : std_logic;
	FA2183 : full_adder port map (N6_1_86,N6_2_86,N6_3_86,N7_2_86,N7_3_87);
-- In matrix 6 adding FA to column 87 
	-- signal N7_0_87 : std_logic;
	-- signal N7_1_88 : std_logic;
	FA2184 : full_adder port map (N5_8_87,N5_9_87,N6_0_87,N7_0_87,N7_1_88);
-- In matrix 6 adding FA to column 87 
	-- signal N7_2_87 : std_logic;
	-- signal N7_3_88 : std_logic;
	FA2185 : full_adder port map (N6_1_87,N6_2_87,N6_3_87,N7_2_87,N7_3_88);
-- In matrix 6 adding FA to column 88 
	-- signal N7_0_88 : std_logic;
	-- signal N7_1_89 : std_logic;
	FA2186 : full_adder port map (N5_8_88,N5_9_88,N6_0_88,N7_0_88,N7_1_89);
-- In matrix 6 adding FA to column 88 
	-- signal N7_2_88 : std_logic;
	-- signal N7_3_89 : std_logic;
	FA2187 : full_adder port map (N6_1_88,N6_2_88,N6_3_88,N7_2_88,N7_3_89);
-- In matrix 6 adding FA to column 89 
	-- signal N7_0_89 : std_logic;
	-- signal N7_1_90 : std_logic;
	FA2188 : full_adder port map (N5_8_89,N5_9_89,N6_0_89,N7_0_89,N7_1_90);
-- In matrix 6 adding FA to column 89 
	-- signal N7_2_89 : std_logic;
	-- signal N7_3_90 : std_logic;
	FA2189 : full_adder port map (N6_1_89,N6_2_89,N6_3_89,N7_2_89,N7_3_90);
-- In matrix 6 adding FA to column 90 
	-- signal N7_0_90 : std_logic;
	-- signal N7_1_91 : std_logic;
	FA2190 : full_adder port map (N5_8_90,N5_9_90,N6_0_90,N7_0_90,N7_1_91);
-- In matrix 6 adding FA to column 90 
	-- signal N7_2_90 : std_logic;
	-- signal N7_3_91 : std_logic;
	FA2191 : full_adder port map (N6_1_90,N6_2_90,N6_3_90,N7_2_90,N7_3_91);
-- In matrix 6 adding FA to column 91 
	-- signal N7_0_91 : std_logic;
	-- signal N7_1_92 : std_logic;
	FA2192 : full_adder port map (N5_7_91,N5_9_91,N6_0_91,N7_0_91,N7_1_92);
-- In matrix 6 adding FA to column 91 
	-- signal N7_2_91 : std_logic;
	-- signal N7_3_92 : std_logic;
	FA2193 : full_adder port map (N6_1_91,N6_2_91,N6_3_91,N7_2_91,N7_3_92);
-- In matrix 6 adding FA to column 92 
	-- signal N7_0_92 : std_logic;
	-- signal N7_1_93 : std_logic;
	FA2194 : full_adder port map (N5_5_92,N5_7_92,N6_0_92,N7_0_92,N7_1_93);
-- In matrix 6 adding FA to column 92 
	-- signal N7_2_92 : std_logic;
	-- signal N7_3_93 : std_logic;
	FA2195 : full_adder port map (N6_1_92,N6_2_92,N6_3_92,N7_2_92,N7_3_93);
-- In matrix 6 adding FA to column 93 
	-- signal N7_0_93 : std_logic;
	-- signal N7_1_94 : std_logic;
	FA2196 : full_adder port map (N5_3_93,N5_5_93,N6_0_93,N7_0_93,N7_1_94);
-- In matrix 6 adding FA to column 93 
	-- signal N7_2_93 : std_logic;
	-- signal N7_3_94 : std_logic;
	FA2197 : full_adder port map (N6_1_93,N6_2_93,N6_3_93,N7_2_93,N7_3_94);
-- In matrix 6 adding FA to column 94 
	-- signal N7_0_94 : std_logic;
	-- signal N7_1_95 : std_logic;
	FA2198 : full_adder port map (N5_1_94,N5_3_94,N6_0_94,N7_0_94,N7_1_95);
-- In matrix 6 adding FA to column 94 
	-- signal N7_2_94 : std_logic;
	-- signal N7_3_95 : std_logic;
	FA2199 : full_adder port map (N6_1_94,N6_2_94,N6_3_94,N7_2_94,N7_3_95);
-- In matrix 6 adding FA to column 95 
	-- signal N7_0_95 : std_logic;
	-- signal N7_1_96 : std_logic;
	FA2200 : full_adder port map (N0_52_95,N5_1_95,N6_0_95,N7_0_95,N7_1_96);
-- In matrix 6 adding FA to column 95 
	-- signal N7_2_95 : std_logic;
	-- signal N7_3_96 : std_logic;
	FA2201 : full_adder port map (N6_1_95,N6_2_95,N6_3_95,N7_2_95,N7_3_96);
-- In matrix 6 adding FA to column 96 
	-- signal N7_0_96 : std_logic;
	-- signal N7_1_97 : std_logic;
	FA2202 : full_adder port map (N0_50_96,N0_51_96,N0_52_96,N7_0_96,N7_1_97);
-- In matrix 6 adding FA to column 96 
	-- signal N7_2_96 : std_logic;
	-- signal N7_3_97 : std_logic;
	FA2203 : full_adder port map (N6_0_96,N6_1_96,N6_2_96,N7_2_96,N7_3_97);
-- In matrix 6 adding FA to column 97 
	-- signal N7_0_97 : std_logic;
	-- signal N7_1_98 : std_logic;
	FA2204 : full_adder port map (N0_48_97,N0_49_97,N0_50_97,N7_0_97,N7_1_98);
-- In matrix 6 adding FA to column 97 
	-- signal N7_2_97 : std_logic;
	-- signal N7_3_98 : std_logic;
	FA2205 : full_adder port map (N0_51_97,N0_52_97,N6_0_97,N7_2_97,N7_3_98);
-- In matrix 6 adding FA to column 98 
	-- signal N7_0_98 : std_logic;
	-- signal N7_1_99 : std_logic;
	FA2206 : full_adder port map (N0_46_98,N0_47_98,N0_48_98,N7_0_98,N7_1_99);
-- In matrix 6 adding FA to column 98 
	-- signal N7_2_98 : std_logic;
	-- signal N7_3_99 : std_logic;
	FA2207 : full_adder port map (N0_49_98,N0_50_98,N0_51_98,N7_2_98,N7_3_99);
-- In matrix 6 adding FA to column 99 
	-- signal N7_0_99 : std_logic;
	-- signal N7_1_100 : std_logic;
	FA2208 : full_adder port map (N0_47_99,N0_48_99,N0_49_99,N7_0_99,N7_1_100);
	-- Elements from matrix 7 
-- In matrix 7 adding HA to column 4 
	-- signal N8_0_4 : std_logic;
	-- signal N8_1_5 : std_logic;
	HA49 : half_adder port map (N0_0_4,N0_1_4,N8_0_4,N8_1_5);
-- In matrix 7 adding FA to column 5 
	-- signal N8_0_5 : std_logic;
	-- signal N8_1_6 : std_logic;
	FA2209 : full_adder port map (N0_0_5,N0_1_5,N0_2_5,N8_0_5,N8_1_6);
-- In matrix 7 adding HA to column 5 
	-- signal N8_2_5 : std_logic;
	-- signal N8_3_6 : std_logic;
	HA50 : half_adder port map (N0_3_5,N0_4_5,N8_2_5,N8_3_6);
-- In matrix 7 adding FA to column 6 
	-- signal N8_0_6 : std_logic;
	-- signal N8_1_7 : std_logic;
	FA2210 : full_adder port map (N0_2_6,N0_3_6,N0_4_6,N8_0_6,N8_1_7);
-- In matrix 7 adding FA to column 6 
	-- signal N8_2_6 : std_logic;
	-- signal N8_3_7 : std_logic;
	FA2211 : full_adder port map (N0_5_6,N0_6_6,N7_0_6,N8_2_6,N8_3_7);
-- In matrix 7 adding FA to column 7 
	-- signal N8_0_7 : std_logic;
	-- signal N8_1_8 : std_logic;
	FA2212 : full_adder port map (N0_5_7,N0_6_7,N0_7_7,N8_0_7,N8_1_8);
-- In matrix 7 adding FA to column 7 
	-- signal N8_2_7 : std_logic;
	-- signal N8_3_8 : std_logic;
	FA2213 : full_adder port map (N7_0_7,N7_1_7,N7_2_7,N8_2_7,N8_3_8);
-- In matrix 7 adding FA to column 8 
	-- signal N8_0_8 : std_logic;
	-- signal N8_1_9 : std_logic;
	FA2214 : full_adder port map (N0_8_8,N6_0_8,N7_0_8,N8_0_8,N8_1_9);
-- In matrix 7 adding FA to column 8 
	-- signal N8_2_8 : std_logic;
	-- signal N8_3_9 : std_logic;
	FA2215 : full_adder port map (N7_1_8,N7_2_8,N7_3_8,N8_2_8,N8_3_9);
-- In matrix 7 adding FA to column 9 
	-- signal N8_0_9 : std_logic;
	-- signal N8_1_10 : std_logic;
	FA2216 : full_adder port map (N6_1_9,N6_2_9,N7_0_9,N8_0_9,N8_1_10);
-- In matrix 7 adding FA to column 9 
	-- signal N8_2_9 : std_logic;
	-- signal N8_3_10 : std_logic;
	FA2217 : full_adder port map (N7_1_9,N7_2_9,N7_3_9,N8_2_9,N8_3_10);
-- In matrix 7 adding FA to column 10 
	-- signal N8_0_10 : std_logic;
	-- signal N8_1_11 : std_logic;
	FA2218 : full_adder port map (N6_3_10,N6_4_10,N7_0_10,N8_0_10,N8_1_11);
-- In matrix 7 adding FA to column 10 
	-- signal N8_2_10 : std_logic;
	-- signal N8_3_11 : std_logic;
	FA2219 : full_adder port map (N7_1_10,N7_2_10,N7_3_10,N8_2_10,N8_3_11);
-- In matrix 7 adding FA to column 11 
	-- signal N8_0_11 : std_logic;
	-- signal N8_1_12 : std_logic;
	FA2220 : full_adder port map (N6_4_11,N6_5_11,N7_0_11,N8_0_11,N8_1_12);
-- In matrix 7 adding FA to column 11 
	-- signal N8_2_11 : std_logic;
	-- signal N8_3_12 : std_logic;
	FA2221 : full_adder port map (N7_1_11,N7_2_11,N7_3_11,N8_2_11,N8_3_12);
-- In matrix 7 adding FA to column 12 
	-- signal N8_0_12 : std_logic;
	-- signal N8_1_13 : std_logic;
	FA2222 : full_adder port map (N6_4_12,N6_5_12,N7_0_12,N8_0_12,N8_1_13);
-- In matrix 7 adding FA to column 12 
	-- signal N8_2_12 : std_logic;
	-- signal N8_3_13 : std_logic;
	FA2223 : full_adder port map (N7_1_12,N7_2_12,N7_3_12,N8_2_12,N8_3_13);
-- In matrix 7 adding FA to column 13 
	-- signal N8_0_13 : std_logic;
	-- signal N8_1_14 : std_logic;
	FA2224 : full_adder port map (N6_4_13,N6_5_13,N7_0_13,N8_0_13,N8_1_14);
-- In matrix 7 adding FA to column 13 
	-- signal N8_2_13 : std_logic;
	-- signal N8_3_14 : std_logic;
	FA2225 : full_adder port map (N7_1_13,N7_2_13,N7_3_13,N8_2_13,N8_3_14);
-- In matrix 7 adding FA to column 14 
	-- signal N8_0_14 : std_logic;
	-- signal N8_1_15 : std_logic;
	FA2226 : full_adder port map (N6_4_14,N6_5_14,N7_0_14,N8_0_14,N8_1_15);
-- In matrix 7 adding FA to column 14 
	-- signal N8_2_14 : std_logic;
	-- signal N8_3_15 : std_logic;
	FA2227 : full_adder port map (N7_1_14,N7_2_14,N7_3_14,N8_2_14,N8_3_15);
-- In matrix 7 adding FA to column 15 
	-- signal N8_0_15 : std_logic;
	-- signal N8_1_16 : std_logic;
	FA2228 : full_adder port map (N6_4_15,N6_5_15,N7_0_15,N8_0_15,N8_1_16);
-- In matrix 7 adding FA to column 15 
	-- signal N8_2_15 : std_logic;
	-- signal N8_3_16 : std_logic;
	FA2229 : full_adder port map (N7_1_15,N7_2_15,N7_3_15,N8_2_15,N8_3_16);
-- In matrix 7 adding FA to column 16 
	-- signal N8_0_16 : std_logic;
	-- signal N8_1_17 : std_logic;
	FA2230 : full_adder port map (N6_4_16,N6_5_16,N7_0_16,N8_0_16,N8_1_17);
-- In matrix 7 adding FA to column 16 
	-- signal N8_2_16 : std_logic;
	-- signal N8_3_17 : std_logic;
	FA2231 : full_adder port map (N7_1_16,N7_2_16,N7_3_16,N8_2_16,N8_3_17);
-- In matrix 7 adding FA to column 17 
	-- signal N8_0_17 : std_logic;
	-- signal N8_1_18 : std_logic;
	FA2232 : full_adder port map (N6_4_17,N6_5_17,N7_0_17,N8_0_17,N8_1_18);
-- In matrix 7 adding FA to column 17 
	-- signal N8_2_17 : std_logic;
	-- signal N8_3_18 : std_logic;
	FA2233 : full_adder port map (N7_1_17,N7_2_17,N7_3_17,N8_2_17,N8_3_18);
-- In matrix 7 adding FA to column 18 
	-- signal N8_0_18 : std_logic;
	-- signal N8_1_19 : std_logic;
	FA2234 : full_adder port map (N6_4_18,N6_5_18,N7_0_18,N8_0_18,N8_1_19);
-- In matrix 7 adding FA to column 18 
	-- signal N8_2_18 : std_logic;
	-- signal N8_3_19 : std_logic;
	FA2235 : full_adder port map (N7_1_18,N7_2_18,N7_3_18,N8_2_18,N8_3_19);
-- In matrix 7 adding FA to column 19 
	-- signal N8_0_19 : std_logic;
	-- signal N8_1_20 : std_logic;
	FA2236 : full_adder port map (N6_4_19,N6_5_19,N7_0_19,N8_0_19,N8_1_20);
-- In matrix 7 adding FA to column 19 
	-- signal N8_2_19 : std_logic;
	-- signal N8_3_20 : std_logic;
	FA2237 : full_adder port map (N7_1_19,N7_2_19,N7_3_19,N8_2_19,N8_3_20);
-- In matrix 7 adding FA to column 20 
	-- signal N8_0_20 : std_logic;
	-- signal N8_1_21 : std_logic;
	FA2238 : full_adder port map (N6_4_20,N6_5_20,N7_0_20,N8_0_20,N8_1_21);
-- In matrix 7 adding FA to column 20 
	-- signal N8_2_20 : std_logic;
	-- signal N8_3_21 : std_logic;
	FA2239 : full_adder port map (N7_1_20,N7_2_20,N7_3_20,N8_2_20,N8_3_21);
-- In matrix 7 adding FA to column 21 
	-- signal N8_0_21 : std_logic;
	-- signal N8_1_22 : std_logic;
	FA2240 : full_adder port map (N6_4_21,N6_5_21,N7_0_21,N8_0_21,N8_1_22);
-- In matrix 7 adding FA to column 21 
	-- signal N8_2_21 : std_logic;
	-- signal N8_3_22 : std_logic;
	FA2241 : full_adder port map (N7_1_21,N7_2_21,N7_3_21,N8_2_21,N8_3_22);
-- In matrix 7 adding FA to column 22 
	-- signal N8_0_22 : std_logic;
	-- signal N8_1_23 : std_logic;
	FA2242 : full_adder port map (N6_4_22,N6_5_22,N7_0_22,N8_0_22,N8_1_23);
-- In matrix 7 adding FA to column 22 
	-- signal N8_2_22 : std_logic;
	-- signal N8_3_23 : std_logic;
	FA2243 : full_adder port map (N7_1_22,N7_2_22,N7_3_22,N8_2_22,N8_3_23);
-- In matrix 7 adding FA to column 23 
	-- signal N8_0_23 : std_logic;
	-- signal N8_1_24 : std_logic;
	FA2244 : full_adder port map (N6_4_23,N6_5_23,N7_0_23,N8_0_23,N8_1_24);
-- In matrix 7 adding FA to column 23 
	-- signal N8_2_23 : std_logic;
	-- signal N8_3_24 : std_logic;
	FA2245 : full_adder port map (N7_1_23,N7_2_23,N7_3_23,N8_2_23,N8_3_24);
-- In matrix 7 adding FA to column 24 
	-- signal N8_0_24 : std_logic;
	-- signal N8_1_25 : std_logic;
	FA2246 : full_adder port map (N6_4_24,N6_5_24,N7_0_24,N8_0_24,N8_1_25);
-- In matrix 7 adding FA to column 24 
	-- signal N8_2_24 : std_logic;
	-- signal N8_3_25 : std_logic;
	FA2247 : full_adder port map (N7_1_24,N7_2_24,N7_3_24,N8_2_24,N8_3_25);
-- In matrix 7 adding FA to column 25 
	-- signal N8_0_25 : std_logic;
	-- signal N8_1_26 : std_logic;
	FA2248 : full_adder port map (N6_4_25,N6_5_25,N7_0_25,N8_0_25,N8_1_26);
-- In matrix 7 adding FA to column 25 
	-- signal N8_2_25 : std_logic;
	-- signal N8_3_26 : std_logic;
	FA2249 : full_adder port map (N7_1_25,N7_2_25,N7_3_25,N8_2_25,N8_3_26);
-- In matrix 7 adding FA to column 26 
	-- signal N8_0_26 : std_logic;
	-- signal N8_1_27 : std_logic;
	FA2250 : full_adder port map (N6_4_26,N6_5_26,N7_0_26,N8_0_26,N8_1_27);
-- In matrix 7 adding FA to column 26 
	-- signal N8_2_26 : std_logic;
	-- signal N8_3_27 : std_logic;
	FA2251 : full_adder port map (N7_1_26,N7_2_26,N7_3_26,N8_2_26,N8_3_27);
-- In matrix 7 adding FA to column 27 
	-- signal N8_0_27 : std_logic;
	-- signal N8_1_28 : std_logic;
	FA2252 : full_adder port map (N6_4_27,N6_5_27,N7_0_27,N8_0_27,N8_1_28);
-- In matrix 7 adding FA to column 27 
	-- signal N8_2_27 : std_logic;
	-- signal N8_3_28 : std_logic;
	FA2253 : full_adder port map (N7_1_27,N7_2_27,N7_3_27,N8_2_27,N8_3_28);
-- In matrix 7 adding FA to column 28 
	-- signal N8_0_28 : std_logic;
	-- signal N8_1_29 : std_logic;
	FA2254 : full_adder port map (N6_4_28,N6_5_28,N7_0_28,N8_0_28,N8_1_29);
-- In matrix 7 adding FA to column 28 
	-- signal N8_2_28 : std_logic;
	-- signal N8_3_29 : std_logic;
	FA2255 : full_adder port map (N7_1_28,N7_2_28,N7_3_28,N8_2_28,N8_3_29);
-- In matrix 7 adding FA to column 29 
	-- signal N8_0_29 : std_logic;
	-- signal N8_1_30 : std_logic;
	FA2256 : full_adder port map (N6_4_29,N6_5_29,N7_0_29,N8_0_29,N8_1_30);
-- In matrix 7 adding FA to column 29 
	-- signal N8_2_29 : std_logic;
	-- signal N8_3_30 : std_logic;
	FA2257 : full_adder port map (N7_1_29,N7_2_29,N7_3_29,N8_2_29,N8_3_30);
-- In matrix 7 adding FA to column 30 
	-- signal N8_0_30 : std_logic;
	-- signal N8_1_31 : std_logic;
	FA2258 : full_adder port map (N6_4_30,N6_5_30,N7_0_30,N8_0_30,N8_1_31);
-- In matrix 7 adding FA to column 30 
	-- signal N8_2_30 : std_logic;
	-- signal N8_3_31 : std_logic;
	FA2259 : full_adder port map (N7_1_30,N7_2_30,N7_3_30,N8_2_30,N8_3_31);
-- In matrix 7 adding FA to column 31 
	-- signal N8_0_31 : std_logic;
	-- signal N8_1_32 : std_logic;
	FA2260 : full_adder port map (N6_4_31,N6_5_31,N7_0_31,N8_0_31,N8_1_32);
-- In matrix 7 adding FA to column 31 
	-- signal N8_2_31 : std_logic;
	-- signal N8_3_32 : std_logic;
	FA2261 : full_adder port map (N7_1_31,N7_2_31,N7_3_31,N8_2_31,N8_3_32);
-- In matrix 7 adding FA to column 32 
	-- signal N8_0_32 : std_logic;
	-- signal N8_1_33 : std_logic;
	FA2262 : full_adder port map (N6_4_32,N6_5_32,N7_0_32,N8_0_32,N8_1_33);
-- In matrix 7 adding FA to column 32 
	-- signal N8_2_32 : std_logic;
	-- signal N8_3_33 : std_logic;
	FA2263 : full_adder port map (N7_1_32,N7_2_32,N7_3_32,N8_2_32,N8_3_33);
-- In matrix 7 adding FA to column 33 
	-- signal N8_0_33 : std_logic;
	-- signal N8_1_34 : std_logic;
	FA2264 : full_adder port map (N6_4_33,N6_5_33,N7_0_33,N8_0_33,N8_1_34);
-- In matrix 7 adding FA to column 33 
	-- signal N8_2_33 : std_logic;
	-- signal N8_3_34 : std_logic;
	FA2265 : full_adder port map (N7_1_33,N7_2_33,N7_3_33,N8_2_33,N8_3_34);
-- In matrix 7 adding FA to column 34 
	-- signal N8_0_34 : std_logic;
	-- signal N8_1_35 : std_logic;
	FA2266 : full_adder port map (N6_4_34,N6_5_34,N7_0_34,N8_0_34,N8_1_35);
-- In matrix 7 adding FA to column 34 
	-- signal N8_2_34 : std_logic;
	-- signal N8_3_35 : std_logic;
	FA2267 : full_adder port map (N7_1_34,N7_2_34,N7_3_34,N8_2_34,N8_3_35);
-- In matrix 7 adding FA to column 35 
	-- signal N8_0_35 : std_logic;
	-- signal N8_1_36 : std_logic;
	FA2268 : full_adder port map (N6_4_35,N6_5_35,N7_0_35,N8_0_35,N8_1_36);
-- In matrix 7 adding FA to column 35 
	-- signal N8_2_35 : std_logic;
	-- signal N8_3_36 : std_logic;
	FA2269 : full_adder port map (N7_1_35,N7_2_35,N7_3_35,N8_2_35,N8_3_36);
-- In matrix 7 adding FA to column 36 
	-- signal N8_0_36 : std_logic;
	-- signal N8_1_37 : std_logic;
	FA2270 : full_adder port map (N6_4_36,N6_5_36,N7_0_36,N8_0_36,N8_1_37);
-- In matrix 7 adding FA to column 36 
	-- signal N8_2_36 : std_logic;
	-- signal N8_3_37 : std_logic;
	FA2271 : full_adder port map (N7_1_36,N7_2_36,N7_3_36,N8_2_36,N8_3_37);
-- In matrix 7 adding FA to column 37 
	-- signal N8_0_37 : std_logic;
	-- signal N8_1_38 : std_logic;
	FA2272 : full_adder port map (N6_4_37,N6_5_37,N7_0_37,N8_0_37,N8_1_38);
-- In matrix 7 adding FA to column 37 
	-- signal N8_2_37 : std_logic;
	-- signal N8_3_38 : std_logic;
	FA2273 : full_adder port map (N7_1_37,N7_2_37,N7_3_37,N8_2_37,N8_3_38);
-- In matrix 7 adding FA to column 38 
	-- signal N8_0_38 : std_logic;
	-- signal N8_1_39 : std_logic;
	FA2274 : full_adder port map (N6_4_38,N6_5_38,N7_0_38,N8_0_38,N8_1_39);
-- In matrix 7 adding FA to column 38 
	-- signal N8_2_38 : std_logic;
	-- signal N8_3_39 : std_logic;
	FA2275 : full_adder port map (N7_1_38,N7_2_38,N7_3_38,N8_2_38,N8_3_39);
-- In matrix 7 adding FA to column 39 
	-- signal N8_0_39 : std_logic;
	-- signal N8_1_40 : std_logic;
	FA2276 : full_adder port map (N6_4_39,N6_5_39,N7_0_39,N8_0_39,N8_1_40);
-- In matrix 7 adding FA to column 39 
	-- signal N8_2_39 : std_logic;
	-- signal N8_3_40 : std_logic;
	FA2277 : full_adder port map (N7_1_39,N7_2_39,N7_3_39,N8_2_39,N8_3_40);
-- In matrix 7 adding FA to column 40 
	-- signal N8_0_40 : std_logic;
	-- signal N8_1_41 : std_logic;
	FA2278 : full_adder port map (N6_4_40,N6_5_40,N7_0_40,N8_0_40,N8_1_41);
-- In matrix 7 adding FA to column 40 
	-- signal N8_2_40 : std_logic;
	-- signal N8_3_41 : std_logic;
	FA2279 : full_adder port map (N7_1_40,N7_2_40,N7_3_40,N8_2_40,N8_3_41);
-- In matrix 7 adding FA to column 41 
	-- signal N8_0_41 : std_logic;
	-- signal N8_1_42 : std_logic;
	FA2280 : full_adder port map (N6_4_41,N6_5_41,N7_0_41,N8_0_41,N8_1_42);
-- In matrix 7 adding FA to column 41 
	-- signal N8_2_41 : std_logic;
	-- signal N8_3_42 : std_logic;
	FA2281 : full_adder port map (N7_1_41,N7_2_41,N7_3_41,N8_2_41,N8_3_42);
-- In matrix 7 adding FA to column 42 
	-- signal N8_0_42 : std_logic;
	-- signal N8_1_43 : std_logic;
	FA2282 : full_adder port map (N6_4_42,N6_5_42,N7_0_42,N8_0_42,N8_1_43);
-- In matrix 7 adding FA to column 42 
	-- signal N8_2_42 : std_logic;
	-- signal N8_3_43 : std_logic;
	FA2283 : full_adder port map (N7_1_42,N7_2_42,N7_3_42,N8_2_42,N8_3_43);
-- In matrix 7 adding FA to column 43 
	-- signal N8_0_43 : std_logic;
	-- signal N8_1_44 : std_logic;
	FA2284 : full_adder port map (N6_4_43,N6_5_43,N7_0_43,N8_0_43,N8_1_44);
-- In matrix 7 adding FA to column 43 
	-- signal N8_2_43 : std_logic;
	-- signal N8_3_44 : std_logic;
	FA2285 : full_adder port map (N7_1_43,N7_2_43,N7_3_43,N8_2_43,N8_3_44);
-- In matrix 7 adding FA to column 44 
	-- signal N8_0_44 : std_logic;
	-- signal N8_1_45 : std_logic;
	FA2286 : full_adder port map (N6_4_44,N6_5_44,N7_0_44,N8_0_44,N8_1_45);
-- In matrix 7 adding FA to column 44 
	-- signal N8_2_44 : std_logic;
	-- signal N8_3_45 : std_logic;
	FA2287 : full_adder port map (N7_1_44,N7_2_44,N7_3_44,N8_2_44,N8_3_45);
-- In matrix 7 adding FA to column 45 
	-- signal N8_0_45 : std_logic;
	-- signal N8_1_46 : std_logic;
	FA2288 : full_adder port map (N6_4_45,N6_5_45,N7_0_45,N8_0_45,N8_1_46);
-- In matrix 7 adding FA to column 45 
	-- signal N8_2_45 : std_logic;
	-- signal N8_3_46 : std_logic;
	FA2289 : full_adder port map (N7_1_45,N7_2_45,N7_3_45,N8_2_45,N8_3_46);
-- In matrix 7 adding FA to column 46 
	-- signal N8_0_46 : std_logic;
	-- signal N8_1_47 : std_logic;
	FA2290 : full_adder port map (N6_4_46,N6_5_46,N7_0_46,N8_0_46,N8_1_47);
-- In matrix 7 adding FA to column 46 
	-- signal N8_2_46 : std_logic;
	-- signal N8_3_47 : std_logic;
	FA2291 : full_adder port map (N7_1_46,N7_2_46,N7_3_46,N8_2_46,N8_3_47);
-- In matrix 7 adding FA to column 47 
	-- signal N8_0_47 : std_logic;
	-- signal N8_1_48 : std_logic;
	FA2292 : full_adder port map (N6_4_47,N6_5_47,N7_0_47,N8_0_47,N8_1_48);
-- In matrix 7 adding FA to column 47 
	-- signal N8_2_47 : std_logic;
	-- signal N8_3_48 : std_logic;
	FA2293 : full_adder port map (N7_1_47,N7_2_47,N7_3_47,N8_2_47,N8_3_48);
-- In matrix 7 adding FA to column 48 
	-- signal N8_0_48 : std_logic;
	-- signal N8_1_49 : std_logic;
	FA2294 : full_adder port map (N6_4_48,N6_5_48,N7_0_48,N8_0_48,N8_1_49);
-- In matrix 7 adding FA to column 48 
	-- signal N8_2_48 : std_logic;
	-- signal N8_3_49 : std_logic;
	FA2295 : full_adder port map (N7_1_48,N7_2_48,N7_3_48,N8_2_48,N8_3_49);
-- In matrix 7 adding FA to column 49 
	-- signal N8_0_49 : std_logic;
	-- signal N8_1_50 : std_logic;
	FA2296 : full_adder port map (N6_4_49,N6_5_49,N7_0_49,N8_0_49,N8_1_50);
-- In matrix 7 adding FA to column 49 
	-- signal N8_2_49 : std_logic;
	-- signal N8_3_50 : std_logic;
	FA2297 : full_adder port map (N7_1_49,N7_2_49,N7_3_49,N8_2_49,N8_3_50);
-- In matrix 7 adding FA to column 50 
	-- signal N8_0_50 : std_logic;
	-- signal N8_1_51 : std_logic;
	FA2298 : full_adder port map (N6_4_50,N6_5_50,N7_0_50,N8_0_50,N8_1_51);
-- In matrix 7 adding FA to column 50 
	-- signal N8_2_50 : std_logic;
	-- signal N8_3_51 : std_logic;
	FA2299 : full_adder port map (N7_1_50,N7_2_50,N7_3_50,N8_2_50,N8_3_51);
-- In matrix 7 adding FA to column 51 
	-- signal N8_0_51 : std_logic;
	-- signal N8_1_52 : std_logic;
	FA2300 : full_adder port map (N6_4_51,N6_5_51,N7_0_51,N8_0_51,N8_1_52);
-- In matrix 7 adding FA to column 51 
	-- signal N8_2_51 : std_logic;
	-- signal N8_3_52 : std_logic;
	FA2301 : full_adder port map (N7_1_51,N7_2_51,N7_3_51,N8_2_51,N8_3_52);
-- In matrix 7 adding FA to column 52 
	-- signal N8_0_52 : std_logic;
	-- signal N8_1_53 : std_logic;
	FA2302 : full_adder port map (N6_4_52,N6_5_52,N7_0_52,N8_0_52,N8_1_53);
-- In matrix 7 adding FA to column 52 
	-- signal N8_2_52 : std_logic;
	-- signal N8_3_53 : std_logic;
	FA2303 : full_adder port map (N7_1_52,N7_2_52,N7_3_52,N8_2_52,N8_3_53);
-- In matrix 7 adding FA to column 53 
	-- signal N8_0_53 : std_logic;
	-- signal N8_1_54 : std_logic;
	FA2304 : full_adder port map (N6_4_53,N6_5_53,N7_0_53,N8_0_53,N8_1_54);
-- In matrix 7 adding FA to column 53 
	-- signal N8_2_53 : std_logic;
	-- signal N8_3_54 : std_logic;
	FA2305 : full_adder port map (N7_1_53,N7_2_53,N7_3_53,N8_2_53,N8_3_54);
-- In matrix 7 adding FA to column 54 
	-- signal N8_0_54 : std_logic;
	-- signal N8_1_55 : std_logic;
	FA2306 : full_adder port map (N6_4_54,N6_5_54,N7_0_54,N8_0_54,N8_1_55);
-- In matrix 7 adding FA to column 54 
	-- signal N8_2_54 : std_logic;
	-- signal N8_3_55 : std_logic;
	FA2307 : full_adder port map (N7_1_54,N7_2_54,N7_3_54,N8_2_54,N8_3_55);
-- In matrix 7 adding FA to column 55 
	-- signal N8_0_55 : std_logic;
	-- signal N8_1_56 : std_logic;
	FA2308 : full_adder port map (N6_4_55,N6_5_55,N7_0_55,N8_0_55,N8_1_56);
-- In matrix 7 adding FA to column 55 
	-- signal N8_2_55 : std_logic;
	-- signal N8_3_56 : std_logic;
	FA2309 : full_adder port map (N7_1_55,N7_2_55,N7_3_55,N8_2_55,N8_3_56);
-- In matrix 7 adding FA to column 56 
	-- signal N8_0_56 : std_logic;
	-- signal N8_1_57 : std_logic;
	FA2310 : full_adder port map (N6_4_56,N6_5_56,N7_0_56,N8_0_56,N8_1_57);
-- In matrix 7 adding FA to column 56 
	-- signal N8_2_56 : std_logic;
	-- signal N8_3_57 : std_logic;
	FA2311 : full_adder port map (N7_1_56,N7_2_56,N7_3_56,N8_2_56,N8_3_57);
-- In matrix 7 adding FA to column 57 
	-- signal N8_0_57 : std_logic;
	-- signal N8_1_58 : std_logic;
	FA2312 : full_adder port map (N6_4_57,N6_5_57,N7_0_57,N8_0_57,N8_1_58);
-- In matrix 7 adding FA to column 57 
	-- signal N8_2_57 : std_logic;
	-- signal N8_3_58 : std_logic;
	FA2313 : full_adder port map (N7_1_57,N7_2_57,N7_3_57,N8_2_57,N8_3_58);
-- In matrix 7 adding FA to column 58 
	-- signal N8_0_58 : std_logic;
	-- signal N8_1_59 : std_logic;
	FA2314 : full_adder port map (N6_4_58,N6_5_58,N7_0_58,N8_0_58,N8_1_59);
-- In matrix 7 adding FA to column 58 
	-- signal N8_2_58 : std_logic;
	-- signal N8_3_59 : std_logic;
	FA2315 : full_adder port map (N7_1_58,N7_2_58,N7_3_58,N8_2_58,N8_3_59);
-- In matrix 7 adding FA to column 59 
	-- signal N8_0_59 : std_logic;
	-- signal N8_1_60 : std_logic;
	FA2316 : full_adder port map (N6_4_59,N6_5_59,N7_0_59,N8_0_59,N8_1_60);
-- In matrix 7 adding FA to column 59 
	-- signal N8_2_59 : std_logic;
	-- signal N8_3_60 : std_logic;
	FA2317 : full_adder port map (N7_1_59,N7_2_59,N7_3_59,N8_2_59,N8_3_60);
-- In matrix 7 adding FA to column 60 
	-- signal N8_0_60 : std_logic;
	-- signal N8_1_61 : std_logic;
	FA2318 : full_adder port map (N6_4_60,N6_5_60,N7_0_60,N8_0_60,N8_1_61);
-- In matrix 7 adding FA to column 60 
	-- signal N8_2_60 : std_logic;
	-- signal N8_3_61 : std_logic;
	FA2319 : full_adder port map (N7_1_60,N7_2_60,N7_3_60,N8_2_60,N8_3_61);
-- In matrix 7 adding FA to column 61 
	-- signal N8_0_61 : std_logic;
	-- signal N8_1_62 : std_logic;
	FA2320 : full_adder port map (N6_4_61,N6_5_61,N7_0_61,N8_0_61,N8_1_62);
-- In matrix 7 adding FA to column 61 
	-- signal N8_2_61 : std_logic;
	-- signal N8_3_62 : std_logic;
	FA2321 : full_adder port map (N7_1_61,N7_2_61,N7_3_61,N8_2_61,N8_3_62);
-- In matrix 7 adding FA to column 62 
	-- signal N8_0_62 : std_logic;
	-- signal N8_1_63 : std_logic;
	FA2322 : full_adder port map (N6_4_62,N6_5_62,N7_0_62,N8_0_62,N8_1_63);
-- In matrix 7 adding FA to column 62 
	-- signal N8_2_62 : std_logic;
	-- signal N8_3_63 : std_logic;
	FA2323 : full_adder port map (N7_1_62,N7_2_62,N7_3_62,N8_2_62,N8_3_63);
-- In matrix 7 adding FA to column 63 
	-- signal N8_0_63 : std_logic;
	-- signal N8_1_64 : std_logic;
	FA2324 : full_adder port map (N6_4_63,N6_5_63,N7_0_63,N8_0_63,N8_1_64);
-- In matrix 7 adding FA to column 63 
	-- signal N8_2_63 : std_logic;
	-- signal N8_3_64 : std_logic;
	FA2325 : full_adder port map (N7_1_63,N7_2_63,N7_3_63,N8_2_63,N8_3_64);
-- In matrix 7 adding FA to column 64 
	-- signal N8_0_64 : std_logic;
	-- signal N8_1_65 : std_logic;
	FA2326 : full_adder port map (N6_4_64,N6_5_64,N7_0_64,N8_0_64,N8_1_65);
-- In matrix 7 adding FA to column 64 
	-- signal N8_2_64 : std_logic;
	-- signal N8_3_65 : std_logic;
	FA2327 : full_adder port map (N7_1_64,N7_2_64,N7_3_64,N8_2_64,N8_3_65);
-- In matrix 7 adding FA to column 65 
	-- signal N8_0_65 : std_logic;
	-- signal N8_1_66 : std_logic;
	FA2328 : full_adder port map (N6_4_65,N6_5_65,N7_0_65,N8_0_65,N8_1_66);
-- In matrix 7 adding FA to column 65 
	-- signal N8_2_65 : std_logic;
	-- signal N8_3_66 : std_logic;
	FA2329 : full_adder port map (N7_1_65,N7_2_65,N7_3_65,N8_2_65,N8_3_66);
-- In matrix 7 adding FA to column 66 
	-- signal N8_0_66 : std_logic;
	-- signal N8_1_67 : std_logic;
	FA2330 : full_adder port map (N6_4_66,N6_5_66,N7_0_66,N8_0_66,N8_1_67);
-- In matrix 7 adding FA to column 66 
	-- signal N8_2_66 : std_logic;
	-- signal N8_3_67 : std_logic;
	FA2331 : full_adder port map (N7_1_66,N7_2_66,N7_3_66,N8_2_66,N8_3_67);
-- In matrix 7 adding FA to column 67 
	-- signal N8_0_67 : std_logic;
	-- signal N8_1_68 : std_logic;
	FA2332 : full_adder port map (N6_4_67,N6_5_67,N7_0_67,N8_0_67,N8_1_68);
-- In matrix 7 adding FA to column 67 
	-- signal N8_2_67 : std_logic;
	-- signal N8_3_68 : std_logic;
	FA2333 : full_adder port map (N7_1_67,N7_2_67,N7_3_67,N8_2_67,N8_3_68);
-- In matrix 7 adding FA to column 68 
	-- signal N8_0_68 : std_logic;
	-- signal N8_1_69 : std_logic;
	FA2334 : full_adder port map (N6_4_68,N6_5_68,N7_0_68,N8_0_68,N8_1_69);
-- In matrix 7 adding FA to column 68 
	-- signal N8_2_68 : std_logic;
	-- signal N8_3_69 : std_logic;
	FA2335 : full_adder port map (N7_1_68,N7_2_68,N7_3_68,N8_2_68,N8_3_69);
-- In matrix 7 adding FA to column 69 
	-- signal N8_0_69 : std_logic;
	-- signal N8_1_70 : std_logic;
	FA2336 : full_adder port map (N6_4_69,N6_5_69,N7_0_69,N8_0_69,N8_1_70);
-- In matrix 7 adding FA to column 69 
	-- signal N8_2_69 : std_logic;
	-- signal N8_3_70 : std_logic;
	FA2337 : full_adder port map (N7_1_69,N7_2_69,N7_3_69,N8_2_69,N8_3_70);
-- In matrix 7 adding FA to column 70 
	-- signal N8_0_70 : std_logic;
	-- signal N8_1_71 : std_logic;
	FA2338 : full_adder port map (N6_4_70,N6_5_70,N7_0_70,N8_0_70,N8_1_71);
-- In matrix 7 adding FA to column 70 
	-- signal N8_2_70 : std_logic;
	-- signal N8_3_71 : std_logic;
	FA2339 : full_adder port map (N7_1_70,N7_2_70,N7_3_70,N8_2_70,N8_3_71);
-- In matrix 7 adding FA to column 71 
	-- signal N8_0_71 : std_logic;
	-- signal N8_1_72 : std_logic;
	FA2340 : full_adder port map (N6_4_71,N6_5_71,N7_0_71,N8_0_71,N8_1_72);
-- In matrix 7 adding FA to column 71 
	-- signal N8_2_71 : std_logic;
	-- signal N8_3_72 : std_logic;
	FA2341 : full_adder port map (N7_1_71,N7_2_71,N7_3_71,N8_2_71,N8_3_72);
-- In matrix 7 adding FA to column 72 
	-- signal N8_0_72 : std_logic;
	-- signal N8_1_73 : std_logic;
	FA2342 : full_adder port map (N6_4_72,N6_5_72,N7_0_72,N8_0_72,N8_1_73);
-- In matrix 7 adding FA to column 72 
	-- signal N8_2_72 : std_logic;
	-- signal N8_3_73 : std_logic;
	FA2343 : full_adder port map (N7_1_72,N7_2_72,N7_3_72,N8_2_72,N8_3_73);
-- In matrix 7 adding FA to column 73 
	-- signal N8_0_73 : std_logic;
	-- signal N8_1_74 : std_logic;
	FA2344 : full_adder port map (N6_4_73,N6_5_73,N7_0_73,N8_0_73,N8_1_74);
-- In matrix 7 adding FA to column 73 
	-- signal N8_2_73 : std_logic;
	-- signal N8_3_74 : std_logic;
	FA2345 : full_adder port map (N7_1_73,N7_2_73,N7_3_73,N8_2_73,N8_3_74);
-- In matrix 7 adding FA to column 74 
	-- signal N8_0_74 : std_logic;
	-- signal N8_1_75 : std_logic;
	FA2346 : full_adder port map (N6_4_74,N6_5_74,N7_0_74,N8_0_74,N8_1_75);
-- In matrix 7 adding FA to column 74 
	-- signal N8_2_74 : std_logic;
	-- signal N8_3_75 : std_logic;
	FA2347 : full_adder port map (N7_1_74,N7_2_74,N7_3_74,N8_2_74,N8_3_75);
-- In matrix 7 adding FA to column 75 
	-- signal N8_0_75 : std_logic;
	-- signal N8_1_76 : std_logic;
	FA2348 : full_adder port map (N6_4_75,N6_5_75,N7_0_75,N8_0_75,N8_1_76);
-- In matrix 7 adding FA to column 75 
	-- signal N8_2_75 : std_logic;
	-- signal N8_3_76 : std_logic;
	FA2349 : full_adder port map (N7_1_75,N7_2_75,N7_3_75,N8_2_75,N8_3_76);
-- In matrix 7 adding FA to column 76 
	-- signal N8_0_76 : std_logic;
	-- signal N8_1_77 : std_logic;
	FA2350 : full_adder port map (N6_4_76,N6_5_76,N7_0_76,N8_0_76,N8_1_77);
-- In matrix 7 adding FA to column 76 
	-- signal N8_2_76 : std_logic;
	-- signal N8_3_77 : std_logic;
	FA2351 : full_adder port map (N7_1_76,N7_2_76,N7_3_76,N8_2_76,N8_3_77);
-- In matrix 7 adding FA to column 77 
	-- signal N8_0_77 : std_logic;
	-- signal N8_1_78 : std_logic;
	FA2352 : full_adder port map (N6_4_77,N6_5_77,N7_0_77,N8_0_77,N8_1_78);
-- In matrix 7 adding FA to column 77 
	-- signal N8_2_77 : std_logic;
	-- signal N8_3_78 : std_logic;
	FA2353 : full_adder port map (N7_1_77,N7_2_77,N7_3_77,N8_2_77,N8_3_78);
-- In matrix 7 adding FA to column 78 
	-- signal N8_0_78 : std_logic;
	-- signal N8_1_79 : std_logic;
	FA2354 : full_adder port map (N6_4_78,N6_5_78,N7_0_78,N8_0_78,N8_1_79);
-- In matrix 7 adding FA to column 78 
	-- signal N8_2_78 : std_logic;
	-- signal N8_3_79 : std_logic;
	FA2355 : full_adder port map (N7_1_78,N7_2_78,N7_3_78,N8_2_78,N8_3_79);
-- In matrix 7 adding FA to column 79 
	-- signal N8_0_79 : std_logic;
	-- signal N8_1_80 : std_logic;
	FA2356 : full_adder port map (N6_4_79,N6_5_79,N7_0_79,N8_0_79,N8_1_80);
-- In matrix 7 adding FA to column 79 
	-- signal N8_2_79 : std_logic;
	-- signal N8_3_80 : std_logic;
	FA2357 : full_adder port map (N7_1_79,N7_2_79,N7_3_79,N8_2_79,N8_3_80);
-- In matrix 7 adding FA to column 80 
	-- signal N8_0_80 : std_logic;
	-- signal N8_1_81 : std_logic;
	FA2358 : full_adder port map (N6_4_80,N6_5_80,N7_0_80,N8_0_80,N8_1_81);
-- In matrix 7 adding FA to column 80 
	-- signal N8_2_80 : std_logic;
	-- signal N8_3_81 : std_logic;
	FA2359 : full_adder port map (N7_1_80,N7_2_80,N7_3_80,N8_2_80,N8_3_81);
-- In matrix 7 adding FA to column 81 
	-- signal N8_0_81 : std_logic;
	-- signal N8_1_82 : std_logic;
	FA2360 : full_adder port map (N6_4_81,N6_5_81,N7_0_81,N8_0_81,N8_1_82);
-- In matrix 7 adding FA to column 81 
	-- signal N8_2_81 : std_logic;
	-- signal N8_3_82 : std_logic;
	FA2361 : full_adder port map (N7_1_81,N7_2_81,N7_3_81,N8_2_81,N8_3_82);
-- In matrix 7 adding FA to column 82 
	-- signal N8_0_82 : std_logic;
	-- signal N8_1_83 : std_logic;
	FA2362 : full_adder port map (N6_4_82,N6_5_82,N7_0_82,N8_0_82,N8_1_83);
-- In matrix 7 adding FA to column 82 
	-- signal N8_2_82 : std_logic;
	-- signal N8_3_83 : std_logic;
	FA2363 : full_adder port map (N7_1_82,N7_2_82,N7_3_82,N8_2_82,N8_3_83);
-- In matrix 7 adding FA to column 83 
	-- signal N8_0_83 : std_logic;
	-- signal N8_1_84 : std_logic;
	FA2364 : full_adder port map (N6_4_83,N6_5_83,N7_0_83,N8_0_83,N8_1_84);
-- In matrix 7 adding FA to column 83 
	-- signal N8_2_83 : std_logic;
	-- signal N8_3_84 : std_logic;
	FA2365 : full_adder port map (N7_1_83,N7_2_83,N7_3_83,N8_2_83,N8_3_84);
-- In matrix 7 adding FA to column 84 
	-- signal N8_0_84 : std_logic;
	-- signal N8_1_85 : std_logic;
	FA2366 : full_adder port map (N6_4_84,N6_5_84,N7_0_84,N8_0_84,N8_1_85);
-- In matrix 7 adding FA to column 84 
	-- signal N8_2_84 : std_logic;
	-- signal N8_3_85 : std_logic;
	FA2367 : full_adder port map (N7_1_84,N7_2_84,N7_3_84,N8_2_84,N8_3_85);
-- In matrix 7 adding FA to column 85 
	-- signal N8_0_85 : std_logic;
	-- signal N8_1_86 : std_logic;
	FA2368 : full_adder port map (N6_4_85,N6_5_85,N7_0_85,N8_0_85,N8_1_86);
-- In matrix 7 adding FA to column 85 
	-- signal N8_2_85 : std_logic;
	-- signal N8_3_86 : std_logic;
	FA2369 : full_adder port map (N7_1_85,N7_2_85,N7_3_85,N8_2_85,N8_3_86);
-- In matrix 7 adding FA to column 86 
	-- signal N8_0_86 : std_logic;
	-- signal N8_1_87 : std_logic;
	FA2370 : full_adder port map (N6_4_86,N6_5_86,N7_0_86,N8_0_86,N8_1_87);
-- In matrix 7 adding FA to column 86 
	-- signal N8_2_86 : std_logic;
	-- signal N8_3_87 : std_logic;
	FA2371 : full_adder port map (N7_1_86,N7_2_86,N7_3_86,N8_2_86,N8_3_87);
-- In matrix 7 adding FA to column 87 
	-- signal N8_0_87 : std_logic;
	-- signal N8_1_88 : std_logic;
	FA2372 : full_adder port map (N6_4_87,N6_5_87,N7_0_87,N8_0_87,N8_1_88);
-- In matrix 7 adding FA to column 87 
	-- signal N8_2_87 : std_logic;
	-- signal N8_3_88 : std_logic;
	FA2373 : full_adder port map (N7_1_87,N7_2_87,N7_3_87,N8_2_87,N8_3_88);
-- In matrix 7 adding FA to column 88 
	-- signal N8_0_88 : std_logic;
	-- signal N8_1_89 : std_logic;
	FA2374 : full_adder port map (N6_4_88,N6_5_88,N7_0_88,N8_0_88,N8_1_89);
-- In matrix 7 adding FA to column 88 
	-- signal N8_2_88 : std_logic;
	-- signal N8_3_89 : std_logic;
	FA2375 : full_adder port map (N7_1_88,N7_2_88,N7_3_88,N8_2_88,N8_3_89);
-- In matrix 7 adding FA to column 89 
	-- signal N8_0_89 : std_logic;
	-- signal N8_1_90 : std_logic;
	FA2376 : full_adder port map (N6_4_89,N6_5_89,N7_0_89,N8_0_89,N8_1_90);
-- In matrix 7 adding FA to column 89 
	-- signal N8_2_89 : std_logic;
	-- signal N8_3_90 : std_logic;
	FA2377 : full_adder port map (N7_1_89,N7_2_89,N7_3_89,N8_2_89,N8_3_90);
-- In matrix 7 adding FA to column 90 
	-- signal N8_0_90 : std_logic;
	-- signal N8_1_91 : std_logic;
	FA2378 : full_adder port map (N6_4_90,N6_5_90,N7_0_90,N8_0_90,N8_1_91);
-- In matrix 7 adding FA to column 90 
	-- signal N8_2_90 : std_logic;
	-- signal N8_3_91 : std_logic;
	FA2379 : full_adder port map (N7_1_90,N7_2_90,N7_3_90,N8_2_90,N8_3_91);
-- In matrix 7 adding FA to column 91 
	-- signal N8_0_91 : std_logic;
	-- signal N8_1_92 : std_logic;
	FA2380 : full_adder port map (N6_4_91,N6_5_91,N7_0_91,N8_0_91,N8_1_92);
-- In matrix 7 adding FA to column 91 
	-- signal N8_2_91 : std_logic;
	-- signal N8_3_92 : std_logic;
	FA2381 : full_adder port map (N7_1_91,N7_2_91,N7_3_91,N8_2_91,N8_3_92);
-- In matrix 7 adding FA to column 92 
	-- signal N8_0_92 : std_logic;
	-- signal N8_1_93 : std_logic;
	FA2382 : full_adder port map (N6_4_92,N6_5_92,N7_0_92,N8_0_92,N8_1_93);
-- In matrix 7 adding FA to column 92 
	-- signal N8_2_92 : std_logic;
	-- signal N8_3_93 : std_logic;
	FA2383 : full_adder port map (N7_1_92,N7_2_92,N7_3_92,N8_2_92,N8_3_93);
-- In matrix 7 adding FA to column 93 
	-- signal N8_0_93 : std_logic;
	-- signal N8_1_94 : std_logic;
	FA2384 : full_adder port map (N6_4_93,N6_5_93,N7_0_93,N8_0_93,N8_1_94);
-- In matrix 7 adding FA to column 93 
	-- signal N8_2_93 : std_logic;
	-- signal N8_3_94 : std_logic;
	FA2385 : full_adder port map (N7_1_93,N7_2_93,N7_3_93,N8_2_93,N8_3_94);
-- In matrix 7 adding FA to column 94 
	-- signal N8_0_94 : std_logic;
	-- signal N8_1_95 : std_logic;
	FA2386 : full_adder port map (N6_4_94,N6_5_94,N7_0_94,N8_0_94,N8_1_95);
-- In matrix 7 adding FA to column 94 
	-- signal N8_2_94 : std_logic;
	-- signal N8_3_95 : std_logic;
	FA2387 : full_adder port map (N7_1_94,N7_2_94,N7_3_94,N8_2_94,N8_3_95);
-- In matrix 7 adding FA to column 95 
	-- signal N8_0_95 : std_logic;
	-- signal N8_1_96 : std_logic;
	FA2388 : full_adder port map (N6_4_95,N6_5_95,N7_0_95,N8_0_95,N8_1_96);
-- In matrix 7 adding FA to column 95 
	-- signal N8_2_95 : std_logic;
	-- signal N8_3_96 : std_logic;
	FA2389 : full_adder port map (N7_1_95,N7_2_95,N7_3_95,N8_2_95,N8_3_96);
-- In matrix 7 adding FA to column 96 
	-- signal N8_0_96 : std_logic;
	-- signal N8_1_97 : std_logic;
	FA2390 : full_adder port map (N6_3_96,N6_5_96,N7_0_96,N8_0_96,N8_1_97);
-- In matrix 7 adding FA to column 96 
	-- signal N8_2_96 : std_logic;
	-- signal N8_3_97 : std_logic;
	FA2391 : full_adder port map (N7_1_96,N7_2_96,N7_3_96,N8_2_96,N8_3_97);
-- In matrix 7 adding FA to column 97 
	-- signal N8_0_97 : std_logic;
	-- signal N8_1_98 : std_logic;
	FA2392 : full_adder port map (N6_1_97,N6_3_97,N7_0_97,N8_0_97,N8_1_98);
-- In matrix 7 adding FA to column 97 
	-- signal N8_2_97 : std_logic;
	-- signal N8_3_98 : std_logic;
	FA2393 : full_adder port map (N7_1_97,N7_2_97,N7_3_97,N8_2_97,N8_3_98);
-- In matrix 7 adding FA to column 98 
	-- signal N8_0_98 : std_logic;
	-- signal N8_1_99 : std_logic;
	FA2394 : full_adder port map (N0_52_98,N6_1_98,N7_0_98,N8_0_98,N8_1_99);
-- In matrix 7 adding FA to column 98 
	-- signal N8_2_98 : std_logic;
	-- signal N8_3_99 : std_logic;
	FA2395 : full_adder port map (N7_1_98,N7_2_98,N7_3_98,N8_2_98,N8_3_99);
-- In matrix 7 adding FA to column 99 
	-- signal N8_0_99 : std_logic;
	-- signal N8_1_100 : std_logic;
	FA2396 : full_adder port map (N0_50_99,N0_51_99,N0_52_99,N8_0_99,N8_1_100);
-- In matrix 7 adding FA to column 99 
	-- signal N8_2_99 : std_logic;
	-- signal N8_3_100 : std_logic;
	FA2397 : full_adder port map (N7_0_99,N7_1_99,N7_3_99,N8_2_99,N8_3_100);
-- In matrix 7 adding FA to column 100 
	-- signal N8_0_100 : std_logic;
	-- signal N8_1_101 : std_logic;
	FA2398 : full_adder port map (N0_48_100,N0_49_100,N0_50_100,N8_0_100,N8_1_101);
-- In matrix 7 adding FA to column 100 
	-- signal N8_2_100 : std_logic;
	-- signal N8_3_101 : std_logic;
	FA2399 : full_adder port map (N0_51_100,N0_52_100,N7_1_100,N8_2_100,N8_3_101);
-- In matrix 7 adding FA to column 101 
	-- signal N8_0_101 : std_logic;
	-- signal N8_1_102 : std_logic;
	FA2400 : full_adder port map (N0_49_101,N0_50_101,N0_51_101,N8_0_101,N8_1_102);
	-- Elements from matrix 8 
-- In matrix 8 adding HA to column 3 
	-- signal N9_0_3 : std_logic;
	-- signal N9_1_4 : std_logic;
	HA51 : half_adder port map (N0_0_3,N0_1_3,N9_0_3,N9_1_4);
-- In matrix 8 adding FA to column 4 
	-- signal N9_0_4 : std_logic;
	-- signal N9_1_5 : std_logic;
	FA2401 : full_adder port map (N0_2_4,N0_3_4,N0_4_4,N9_0_4,N9_1_5);
-- In matrix 8 adding FA to column 5 
	-- signal N9_0_5 : std_logic;
	-- signal N9_1_6 : std_logic;
	FA2402 : full_adder port map (N0_5_5,N8_0_5,N8_1_5,N9_0_5,N9_1_6);
-- In matrix 8 adding FA to column 6 
	-- signal N9_0_6 : std_logic;
	-- signal N9_1_7 : std_logic;
	FA2403 : full_adder port map (N8_0_6,N8_1_6,N8_2_6,N9_0_6,N9_1_7);
-- In matrix 8 adding FA to column 7 
	-- signal N9_0_7 : std_logic;
	-- signal N9_1_8 : std_logic;
	FA2404 : full_adder port map (N8_0_7,N8_1_7,N8_2_7,N9_0_7,N9_1_8);
-- In matrix 8 adding FA to column 8 
	-- signal N9_0_8 : std_logic;
	-- signal N9_1_9 : std_logic;
	FA2405 : full_adder port map (N8_0_8,N8_1_8,N8_2_8,N9_0_8,N9_1_9);
-- In matrix 8 adding FA to column 9 
	-- signal N9_0_9 : std_logic;
	-- signal N9_1_10 : std_logic;
	FA2406 : full_adder port map (N8_0_9,N8_1_9,N8_2_9,N9_0_9,N9_1_10);
-- In matrix 8 adding FA to column 10 
	-- signal N9_0_10 : std_logic;
	-- signal N9_1_11 : std_logic;
	FA2407 : full_adder port map (N8_0_10,N8_1_10,N8_2_10,N9_0_10,N9_1_11);
-- In matrix 8 adding FA to column 11 
	-- signal N9_0_11 : std_logic;
	-- signal N9_1_12 : std_logic;
	FA2408 : full_adder port map (N8_0_11,N8_1_11,N8_2_11,N9_0_11,N9_1_12);
-- In matrix 8 adding FA to column 12 
	-- signal N9_0_12 : std_logic;
	-- signal N9_1_13 : std_logic;
	FA2409 : full_adder port map (N8_0_12,N8_1_12,N8_2_12,N9_0_12,N9_1_13);
-- In matrix 8 adding FA to column 13 
	-- signal N9_0_13 : std_logic;
	-- signal N9_1_14 : std_logic;
	FA2410 : full_adder port map (N8_0_13,N8_1_13,N8_2_13,N9_0_13,N9_1_14);
-- In matrix 8 adding FA to column 14 
	-- signal N9_0_14 : std_logic;
	-- signal N9_1_15 : std_logic;
	FA2411 : full_adder port map (N8_0_14,N8_1_14,N8_2_14,N9_0_14,N9_1_15);
-- In matrix 8 adding FA to column 15 
	-- signal N9_0_15 : std_logic;
	-- signal N9_1_16 : std_logic;
	FA2412 : full_adder port map (N8_0_15,N8_1_15,N8_2_15,N9_0_15,N9_1_16);
-- In matrix 8 adding FA to column 16 
	-- signal N9_0_16 : std_logic;
	-- signal N9_1_17 : std_logic;
	FA2413 : full_adder port map (N8_0_16,N8_1_16,N8_2_16,N9_0_16,N9_1_17);
-- In matrix 8 adding FA to column 17 
	-- signal N9_0_17 : std_logic;
	-- signal N9_1_18 : std_logic;
	FA2414 : full_adder port map (N8_0_17,N8_1_17,N8_2_17,N9_0_17,N9_1_18);
-- In matrix 8 adding FA to column 18 
	-- signal N9_0_18 : std_logic;
	-- signal N9_1_19 : std_logic;
	FA2415 : full_adder port map (N8_0_18,N8_1_18,N8_2_18,N9_0_18,N9_1_19);
-- In matrix 8 adding FA to column 19 
	-- signal N9_0_19 : std_logic;
	-- signal N9_1_20 : std_logic;
	FA2416 : full_adder port map (N8_0_19,N8_1_19,N8_2_19,N9_0_19,N9_1_20);
-- In matrix 8 adding FA to column 20 
	-- signal N9_0_20 : std_logic;
	-- signal N9_1_21 : std_logic;
	FA2417 : full_adder port map (N8_0_20,N8_1_20,N8_2_20,N9_0_20,N9_1_21);
-- In matrix 8 adding FA to column 21 
	-- signal N9_0_21 : std_logic;
	-- signal N9_1_22 : std_logic;
	FA2418 : full_adder port map (N8_0_21,N8_1_21,N8_2_21,N9_0_21,N9_1_22);
-- In matrix 8 adding FA to column 22 
	-- signal N9_0_22 : std_logic;
	-- signal N9_1_23 : std_logic;
	FA2419 : full_adder port map (N8_0_22,N8_1_22,N8_2_22,N9_0_22,N9_1_23);
-- In matrix 8 adding FA to column 23 
	-- signal N9_0_23 : std_logic;
	-- signal N9_1_24 : std_logic;
	FA2420 : full_adder port map (N8_0_23,N8_1_23,N8_2_23,N9_0_23,N9_1_24);
-- In matrix 8 adding FA to column 24 
	-- signal N9_0_24 : std_logic;
	-- signal N9_1_25 : std_logic;
	FA2421 : full_adder port map (N8_0_24,N8_1_24,N8_2_24,N9_0_24,N9_1_25);
-- In matrix 8 adding FA to column 25 
	-- signal N9_0_25 : std_logic;
	-- signal N9_1_26 : std_logic;
	FA2422 : full_adder port map (N8_0_25,N8_1_25,N8_2_25,N9_0_25,N9_1_26);
-- In matrix 8 adding FA to column 26 
	-- signal N9_0_26 : std_logic;
	-- signal N9_1_27 : std_logic;
	FA2423 : full_adder port map (N8_0_26,N8_1_26,N8_2_26,N9_0_26,N9_1_27);
-- In matrix 8 adding FA to column 27 
	-- signal N9_0_27 : std_logic;
	-- signal N9_1_28 : std_logic;
	FA2424 : full_adder port map (N8_0_27,N8_1_27,N8_2_27,N9_0_27,N9_1_28);
-- In matrix 8 adding FA to column 28 
	-- signal N9_0_28 : std_logic;
	-- signal N9_1_29 : std_logic;
	FA2425 : full_adder port map (N8_0_28,N8_1_28,N8_2_28,N9_0_28,N9_1_29);
-- In matrix 8 adding FA to column 29 
	-- signal N9_0_29 : std_logic;
	-- signal N9_1_30 : std_logic;
	FA2426 : full_adder port map (N8_0_29,N8_1_29,N8_2_29,N9_0_29,N9_1_30);
-- In matrix 8 adding FA to column 30 
	-- signal N9_0_30 : std_logic;
	-- signal N9_1_31 : std_logic;
	FA2427 : full_adder port map (N8_0_30,N8_1_30,N8_2_30,N9_0_30,N9_1_31);
-- In matrix 8 adding FA to column 31 
	-- signal N9_0_31 : std_logic;
	-- signal N9_1_32 : std_logic;
	FA2428 : full_adder port map (N8_0_31,N8_1_31,N8_2_31,N9_0_31,N9_1_32);
-- In matrix 8 adding FA to column 32 
	-- signal N9_0_32 : std_logic;
	-- signal N9_1_33 : std_logic;
	FA2429 : full_adder port map (N8_0_32,N8_1_32,N8_2_32,N9_0_32,N9_1_33);
-- In matrix 8 adding FA to column 33 
	-- signal N9_0_33 : std_logic;
	-- signal N9_1_34 : std_logic;
	FA2430 : full_adder port map (N8_0_33,N8_1_33,N8_2_33,N9_0_33,N9_1_34);
-- In matrix 8 adding FA to column 34 
	-- signal N9_0_34 : std_logic;
	-- signal N9_1_35 : std_logic;
	FA2431 : full_adder port map (N8_0_34,N8_1_34,N8_2_34,N9_0_34,N9_1_35);
-- In matrix 8 adding FA to column 35 
	-- signal N9_0_35 : std_logic;
	-- signal N9_1_36 : std_logic;
	FA2432 : full_adder port map (N8_0_35,N8_1_35,N8_2_35,N9_0_35,N9_1_36);
-- In matrix 8 adding FA to column 36 
	-- signal N9_0_36 : std_logic;
	-- signal N9_1_37 : std_logic;
	FA2433 : full_adder port map (N8_0_36,N8_1_36,N8_2_36,N9_0_36,N9_1_37);
-- In matrix 8 adding FA to column 37 
	-- signal N9_0_37 : std_logic;
	-- signal N9_1_38 : std_logic;
	FA2434 : full_adder port map (N8_0_37,N8_1_37,N8_2_37,N9_0_37,N9_1_38);
-- In matrix 8 adding FA to column 38 
	-- signal N9_0_38 : std_logic;
	-- signal N9_1_39 : std_logic;
	FA2435 : full_adder port map (N8_0_38,N8_1_38,N8_2_38,N9_0_38,N9_1_39);
-- In matrix 8 adding FA to column 39 
	-- signal N9_0_39 : std_logic;
	-- signal N9_1_40 : std_logic;
	FA2436 : full_adder port map (N8_0_39,N8_1_39,N8_2_39,N9_0_39,N9_1_40);
-- In matrix 8 adding FA to column 40 
	-- signal N9_0_40 : std_logic;
	-- signal N9_1_41 : std_logic;
	FA2437 : full_adder port map (N8_0_40,N8_1_40,N8_2_40,N9_0_40,N9_1_41);
-- In matrix 8 adding FA to column 41 
	-- signal N9_0_41 : std_logic;
	-- signal N9_1_42 : std_logic;
	FA2438 : full_adder port map (N8_0_41,N8_1_41,N8_2_41,N9_0_41,N9_1_42);
-- In matrix 8 adding FA to column 42 
	-- signal N9_0_42 : std_logic;
	-- signal N9_1_43 : std_logic;
	FA2439 : full_adder port map (N8_0_42,N8_1_42,N8_2_42,N9_0_42,N9_1_43);
-- In matrix 8 adding FA to column 43 
	-- signal N9_0_43 : std_logic;
	-- signal N9_1_44 : std_logic;
	FA2440 : full_adder port map (N8_0_43,N8_1_43,N8_2_43,N9_0_43,N9_1_44);
-- In matrix 8 adding FA to column 44 
	-- signal N9_0_44 : std_logic;
	-- signal N9_1_45 : std_logic;
	FA2441 : full_adder port map (N8_0_44,N8_1_44,N8_2_44,N9_0_44,N9_1_45);
-- In matrix 8 adding FA to column 45 
	-- signal N9_0_45 : std_logic;
	-- signal N9_1_46 : std_logic;
	FA2442 : full_adder port map (N8_0_45,N8_1_45,N8_2_45,N9_0_45,N9_1_46);
-- In matrix 8 adding FA to column 46 
	-- signal N9_0_46 : std_logic;
	-- signal N9_1_47 : std_logic;
	FA2443 : full_adder port map (N8_0_46,N8_1_46,N8_2_46,N9_0_46,N9_1_47);
-- In matrix 8 adding FA to column 47 
	-- signal N9_0_47 : std_logic;
	-- signal N9_1_48 : std_logic;
	FA2444 : full_adder port map (N8_0_47,N8_1_47,N8_2_47,N9_0_47,N9_1_48);
-- In matrix 8 adding FA to column 48 
	-- signal N9_0_48 : std_logic;
	-- signal N9_1_49 : std_logic;
	FA2445 : full_adder port map (N8_0_48,N8_1_48,N8_2_48,N9_0_48,N9_1_49);
-- In matrix 8 adding FA to column 49 
	-- signal N9_0_49 : std_logic;
	-- signal N9_1_50 : std_logic;
	FA2446 : full_adder port map (N8_0_49,N8_1_49,N8_2_49,N9_0_49,N9_1_50);
-- In matrix 8 adding FA to column 50 
	-- signal N9_0_50 : std_logic;
	-- signal N9_1_51 : std_logic;
	FA2447 : full_adder port map (N8_0_50,N8_1_50,N8_2_50,N9_0_50,N9_1_51);
-- In matrix 8 adding FA to column 51 
	-- signal N9_0_51 : std_logic;
	-- signal N9_1_52 : std_logic;
	FA2448 : full_adder port map (N8_0_51,N8_1_51,N8_2_51,N9_0_51,N9_1_52);
-- In matrix 8 adding FA to column 52 
	-- signal N9_0_52 : std_logic;
	-- signal N9_1_53 : std_logic;
	FA2449 : full_adder port map (N8_0_52,N8_1_52,N8_2_52,N9_0_52,N9_1_53);
-- In matrix 8 adding FA to column 53 
	-- signal N9_0_53 : std_logic;
	-- signal N9_1_54 : std_logic;
	FA2450 : full_adder port map (N8_0_53,N8_1_53,N8_2_53,N9_0_53,N9_1_54);
-- In matrix 8 adding FA to column 54 
	-- signal N9_0_54 : std_logic;
	-- signal N9_1_55 : std_logic;
	FA2451 : full_adder port map (N8_0_54,N8_1_54,N8_2_54,N9_0_54,N9_1_55);
-- In matrix 8 adding FA to column 55 
	-- signal N9_0_55 : std_logic;
	-- signal N9_1_56 : std_logic;
	FA2452 : full_adder port map (N8_0_55,N8_1_55,N8_2_55,N9_0_55,N9_1_56);
-- In matrix 8 adding FA to column 56 
	-- signal N9_0_56 : std_logic;
	-- signal N9_1_57 : std_logic;
	FA2453 : full_adder port map (N8_0_56,N8_1_56,N8_2_56,N9_0_56,N9_1_57);
-- In matrix 8 adding FA to column 57 
	-- signal N9_0_57 : std_logic;
	-- signal N9_1_58 : std_logic;
	FA2454 : full_adder port map (N8_0_57,N8_1_57,N8_2_57,N9_0_57,N9_1_58);
-- In matrix 8 adding FA to column 58 
	-- signal N9_0_58 : std_logic;
	-- signal N9_1_59 : std_logic;
	FA2455 : full_adder port map (N8_0_58,N8_1_58,N8_2_58,N9_0_58,N9_1_59);
-- In matrix 8 adding FA to column 59 
	-- signal N9_0_59 : std_logic;
	-- signal N9_1_60 : std_logic;
	FA2456 : full_adder port map (N8_0_59,N8_1_59,N8_2_59,N9_0_59,N9_1_60);
-- In matrix 8 adding FA to column 60 
	-- signal N9_0_60 : std_logic;
	-- signal N9_1_61 : std_logic;
	FA2457 : full_adder port map (N8_0_60,N8_1_60,N8_2_60,N9_0_60,N9_1_61);
-- In matrix 8 adding FA to column 61 
	-- signal N9_0_61 : std_logic;
	-- signal N9_1_62 : std_logic;
	FA2458 : full_adder port map (N8_0_61,N8_1_61,N8_2_61,N9_0_61,N9_1_62);
-- In matrix 8 adding FA to column 62 
	-- signal N9_0_62 : std_logic;
	-- signal N9_1_63 : std_logic;
	FA2459 : full_adder port map (N8_0_62,N8_1_62,N8_2_62,N9_0_62,N9_1_63);
-- In matrix 8 adding FA to column 63 
	-- signal N9_0_63 : std_logic;
	-- signal N9_1_64 : std_logic;
	FA2460 : full_adder port map (N8_0_63,N8_1_63,N8_2_63,N9_0_63,N9_1_64);
-- In matrix 8 adding FA to column 64 
	-- signal N9_0_64 : std_logic;
	-- signal N9_1_65 : std_logic;
	FA2461 : full_adder port map (N8_0_64,N8_1_64,N8_2_64,N9_0_64,N9_1_65);
-- In matrix 8 adding FA to column 65 
	-- signal N9_0_65 : std_logic;
	-- signal N9_1_66 : std_logic;
	FA2462 : full_adder port map (N8_0_65,N8_1_65,N8_2_65,N9_0_65,N9_1_66);
-- In matrix 8 adding FA to column 66 
	-- signal N9_0_66 : std_logic;
	-- signal N9_1_67 : std_logic;
	FA2463 : full_adder port map (N8_0_66,N8_1_66,N8_2_66,N9_0_66,N9_1_67);
-- In matrix 8 adding FA to column 67 
	-- signal N9_0_67 : std_logic;
	-- signal N9_1_68 : std_logic;
	FA2464 : full_adder port map (N8_0_67,N8_1_67,N8_2_67,N9_0_67,N9_1_68);
-- In matrix 8 adding FA to column 68 
	-- signal N9_0_68 : std_logic;
	-- signal N9_1_69 : std_logic;
	FA2465 : full_adder port map (N8_0_68,N8_1_68,N8_2_68,N9_0_68,N9_1_69);
-- In matrix 8 adding FA to column 69 
	-- signal N9_0_69 : std_logic;
	-- signal N9_1_70 : std_logic;
	FA2466 : full_adder port map (N8_0_69,N8_1_69,N8_2_69,N9_0_69,N9_1_70);
-- In matrix 8 adding FA to column 70 
	-- signal N9_0_70 : std_logic;
	-- signal N9_1_71 : std_logic;
	FA2467 : full_adder port map (N8_0_70,N8_1_70,N8_2_70,N9_0_70,N9_1_71);
-- In matrix 8 adding FA to column 71 
	-- signal N9_0_71 : std_logic;
	-- signal N9_1_72 : std_logic;
	FA2468 : full_adder port map (N8_0_71,N8_1_71,N8_2_71,N9_0_71,N9_1_72);
-- In matrix 8 adding FA to column 72 
	-- signal N9_0_72 : std_logic;
	-- signal N9_1_73 : std_logic;
	FA2469 : full_adder port map (N8_0_72,N8_1_72,N8_2_72,N9_0_72,N9_1_73);
-- In matrix 8 adding FA to column 73 
	-- signal N9_0_73 : std_logic;
	-- signal N9_1_74 : std_logic;
	FA2470 : full_adder port map (N8_0_73,N8_1_73,N8_2_73,N9_0_73,N9_1_74);
-- In matrix 8 adding FA to column 74 
	-- signal N9_0_74 : std_logic;
	-- signal N9_1_75 : std_logic;
	FA2471 : full_adder port map (N8_0_74,N8_1_74,N8_2_74,N9_0_74,N9_1_75);
-- In matrix 8 adding FA to column 75 
	-- signal N9_0_75 : std_logic;
	-- signal N9_1_76 : std_logic;
	FA2472 : full_adder port map (N8_0_75,N8_1_75,N8_2_75,N9_0_75,N9_1_76);
-- In matrix 8 adding FA to column 76 
	-- signal N9_0_76 : std_logic;
	-- signal N9_1_77 : std_logic;
	FA2473 : full_adder port map (N8_0_76,N8_1_76,N8_2_76,N9_0_76,N9_1_77);
-- In matrix 8 adding FA to column 77 
	-- signal N9_0_77 : std_logic;
	-- signal N9_1_78 : std_logic;
	FA2474 : full_adder port map (N8_0_77,N8_1_77,N8_2_77,N9_0_77,N9_1_78);
-- In matrix 8 adding FA to column 78 
	-- signal N9_0_78 : std_logic;
	-- signal N9_1_79 : std_logic;
	FA2475 : full_adder port map (N8_0_78,N8_1_78,N8_2_78,N9_0_78,N9_1_79);
-- In matrix 8 adding FA to column 79 
	-- signal N9_0_79 : std_logic;
	-- signal N9_1_80 : std_logic;
	FA2476 : full_adder port map (N8_0_79,N8_1_79,N8_2_79,N9_0_79,N9_1_80);
-- In matrix 8 adding FA to column 80 
	-- signal N9_0_80 : std_logic;
	-- signal N9_1_81 : std_logic;
	FA2477 : full_adder port map (N8_0_80,N8_1_80,N8_2_80,N9_0_80,N9_1_81);
-- In matrix 8 adding FA to column 81 
	-- signal N9_0_81 : std_logic;
	-- signal N9_1_82 : std_logic;
	FA2478 : full_adder port map (N8_0_81,N8_1_81,N8_2_81,N9_0_81,N9_1_82);
-- In matrix 8 adding FA to column 82 
	-- signal N9_0_82 : std_logic;
	-- signal N9_1_83 : std_logic;
	FA2479 : full_adder port map (N8_0_82,N8_1_82,N8_2_82,N9_0_82,N9_1_83);
-- In matrix 8 adding FA to column 83 
	-- signal N9_0_83 : std_logic;
	-- signal N9_1_84 : std_logic;
	FA2480 : full_adder port map (N8_0_83,N8_1_83,N8_2_83,N9_0_83,N9_1_84);
-- In matrix 8 adding FA to column 84 
	-- signal N9_0_84 : std_logic;
	-- signal N9_1_85 : std_logic;
	FA2481 : full_adder port map (N8_0_84,N8_1_84,N8_2_84,N9_0_84,N9_1_85);
-- In matrix 8 adding FA to column 85 
	-- signal N9_0_85 : std_logic;
	-- signal N9_1_86 : std_logic;
	FA2482 : full_adder port map (N8_0_85,N8_1_85,N8_2_85,N9_0_85,N9_1_86);
-- In matrix 8 adding FA to column 86 
	-- signal N9_0_86 : std_logic;
	-- signal N9_1_87 : std_logic;
	FA2483 : full_adder port map (N8_0_86,N8_1_86,N8_2_86,N9_0_86,N9_1_87);
-- In matrix 8 adding FA to column 87 
	-- signal N9_0_87 : std_logic;
	-- signal N9_1_88 : std_logic;
	FA2484 : full_adder port map (N8_0_87,N8_1_87,N8_2_87,N9_0_87,N9_1_88);
-- In matrix 8 adding FA to column 88 
	-- signal N9_0_88 : std_logic;
	-- signal N9_1_89 : std_logic;
	FA2485 : full_adder port map (N8_0_88,N8_1_88,N8_2_88,N9_0_88,N9_1_89);
-- In matrix 8 adding FA to column 89 
	-- signal N9_0_89 : std_logic;
	-- signal N9_1_90 : std_logic;
	FA2486 : full_adder port map (N8_0_89,N8_1_89,N8_2_89,N9_0_89,N9_1_90);
-- In matrix 8 adding FA to column 90 
	-- signal N9_0_90 : std_logic;
	-- signal N9_1_91 : std_logic;
	FA2487 : full_adder port map (N8_0_90,N8_1_90,N8_2_90,N9_0_90,N9_1_91);
-- In matrix 8 adding FA to column 91 
	-- signal N9_0_91 : std_logic;
	-- signal N9_1_92 : std_logic;
	FA2488 : full_adder port map (N8_0_91,N8_1_91,N8_2_91,N9_0_91,N9_1_92);
-- In matrix 8 adding FA to column 92 
	-- signal N9_0_92 : std_logic;
	-- signal N9_1_93 : std_logic;
	FA2489 : full_adder port map (N8_0_92,N8_1_92,N8_2_92,N9_0_92,N9_1_93);
-- In matrix 8 adding FA to column 93 
	-- signal N9_0_93 : std_logic;
	-- signal N9_1_94 : std_logic;
	FA2490 : full_adder port map (N8_0_93,N8_1_93,N8_2_93,N9_0_93,N9_1_94);
-- In matrix 8 adding FA to column 94 
	-- signal N9_0_94 : std_logic;
	-- signal N9_1_95 : std_logic;
	FA2491 : full_adder port map (N8_0_94,N8_1_94,N8_2_94,N9_0_94,N9_1_95);
-- In matrix 8 adding FA to column 95 
	-- signal N9_0_95 : std_logic;
	-- signal N9_1_96 : std_logic;
	FA2492 : full_adder port map (N8_0_95,N8_1_95,N8_2_95,N9_0_95,N9_1_96);
-- In matrix 8 adding FA to column 96 
	-- signal N9_0_96 : std_logic;
	-- signal N9_1_97 : std_logic;
	FA2493 : full_adder port map (N8_0_96,N8_1_96,N8_2_96,N9_0_96,N9_1_97);
-- In matrix 8 adding FA to column 97 
	-- signal N9_0_97 : std_logic;
	-- signal N9_1_98 : std_logic;
	FA2494 : full_adder port map (N8_0_97,N8_1_97,N8_2_97,N9_0_97,N9_1_98);
-- In matrix 8 adding FA to column 98 
	-- signal N9_0_98 : std_logic;
	-- signal N9_1_99 : std_logic;
	FA2495 : full_adder port map (N8_0_98,N8_1_98,N8_2_98,N9_0_98,N9_1_99);
-- In matrix 8 adding FA to column 99 
	-- signal N9_0_99 : std_logic;
	-- signal N9_1_100 : std_logic;
	FA2496 : full_adder port map (N8_0_99,N8_1_99,N8_2_99,N9_0_99,N9_1_100);
-- In matrix 8 adding FA to column 100 
	-- signal N9_0_100 : std_logic;
	-- signal N9_1_101 : std_logic;
	FA2497 : full_adder port map (N8_0_100,N8_1_100,N8_2_100,N9_0_100,N9_1_101);
-- In matrix 8 adding FA to column 101 
	-- signal N9_0_101 : std_logic;
	-- signal N9_1_102 : std_logic;
	FA2498 : full_adder port map (N0_52_101,N8_0_101,N8_1_101,N9_0_101,N9_1_102);
-- In matrix 8 adding FA to column 102 
	-- signal N9_0_102 : std_logic;
	-- signal N9_1_103 : std_logic;
	FA2499 : full_adder port map (N0_50_102,N0_51_102,N0_52_102,N9_0_102,N9_1_103);
	-- Elements from matrix 9 
-- In matrix 9 adding HA to column 2 
	-- signal N10_0_2 : std_logic;
	-- signal N10_1_3 : std_logic;
	HA52 : half_adder port map (N0_0_2,N0_1_2,N10_0_2,N10_1_3);
-- In matrix 9 adding FA to column 3 
	-- signal N10_0_3 : std_logic;
	-- signal N10_1_4 : std_logic;
	FA2500 : full_adder port map (N0_2_3,N0_3_3,N9_0_3,N10_0_3,N10_1_4);
-- In matrix 9 adding FA to column 4 
	-- signal N10_0_4 : std_logic;
	-- signal N10_1_5 : std_logic;
	FA2501 : full_adder port map (N8_0_4,N9_0_4,N9_1_4,N10_0_4,N10_1_5);
-- In matrix 9 adding FA to column 5 
	-- signal N10_0_5 : std_logic;
	-- signal N10_1_6 : std_logic;
	FA2502 : full_adder port map (N8_2_5,N9_0_5,N9_1_5,N10_0_5,N10_1_6);
-- In matrix 9 adding FA to column 6 
	-- signal N10_0_6 : std_logic;
	-- signal N10_1_7 : std_logic;
	FA2503 : full_adder port map (N8_3_6,N9_0_6,N9_1_6,N10_0_6,N10_1_7);
-- In matrix 9 adding FA to column 7 
	-- signal N10_0_7 : std_logic;
	-- signal N10_1_8 : std_logic;
	FA2504 : full_adder port map (N8_3_7,N9_0_7,N9_1_7,N10_0_7,N10_1_8);
-- In matrix 9 adding FA to column 8 
	-- signal N10_0_8 : std_logic;
	-- signal N10_1_9 : std_logic;
	FA2505 : full_adder port map (N8_3_8,N9_0_8,N9_1_8,N10_0_8,N10_1_9);
-- In matrix 9 adding FA to column 9 
	-- signal N10_0_9 : std_logic;
	-- signal N10_1_10 : std_logic;
	FA2506 : full_adder port map (N8_3_9,N9_0_9,N9_1_9,N10_0_9,N10_1_10);
-- In matrix 9 adding FA to column 10 
	-- signal N10_0_10 : std_logic;
	-- signal N10_1_11 : std_logic;
	FA2507 : full_adder port map (N8_3_10,N9_0_10,N9_1_10,N10_0_10,N10_1_11);
-- In matrix 9 adding FA to column 11 
	-- signal N10_0_11 : std_logic;
	-- signal N10_1_12 : std_logic;
	FA2508 : full_adder port map (N8_3_11,N9_0_11,N9_1_11,N10_0_11,N10_1_12);
-- In matrix 9 adding FA to column 12 
	-- signal N10_0_12 : std_logic;
	-- signal N10_1_13 : std_logic;
	FA2509 : full_adder port map (N8_3_12,N9_0_12,N9_1_12,N10_0_12,N10_1_13);
-- In matrix 9 adding FA to column 13 
	-- signal N10_0_13 : std_logic;
	-- signal N10_1_14 : std_logic;
	FA2510 : full_adder port map (N8_3_13,N9_0_13,N9_1_13,N10_0_13,N10_1_14);
-- In matrix 9 adding FA to column 14 
	-- signal N10_0_14 : std_logic;
	-- signal N10_1_15 : std_logic;
	FA2511 : full_adder port map (N8_3_14,N9_0_14,N9_1_14,N10_0_14,N10_1_15);
-- In matrix 9 adding FA to column 15 
	-- signal N10_0_15 : std_logic;
	-- signal N10_1_16 : std_logic;
	FA2512 : full_adder port map (N8_3_15,N9_0_15,N9_1_15,N10_0_15,N10_1_16);
-- In matrix 9 adding FA to column 16 
	-- signal N10_0_16 : std_logic;
	-- signal N10_1_17 : std_logic;
	FA2513 : full_adder port map (N8_3_16,N9_0_16,N9_1_16,N10_0_16,N10_1_17);
-- In matrix 9 adding FA to column 17 
	-- signal N10_0_17 : std_logic;
	-- signal N10_1_18 : std_logic;
	FA2514 : full_adder port map (N8_3_17,N9_0_17,N9_1_17,N10_0_17,N10_1_18);
-- In matrix 9 adding FA to column 18 
	-- signal N10_0_18 : std_logic;
	-- signal N10_1_19 : std_logic;
	FA2515 : full_adder port map (N8_3_18,N9_0_18,N9_1_18,N10_0_18,N10_1_19);
-- In matrix 9 adding FA to column 19 
	-- signal N10_0_19 : std_logic;
	-- signal N10_1_20 : std_logic;
	FA2516 : full_adder port map (N8_3_19,N9_0_19,N9_1_19,N10_0_19,N10_1_20);
-- In matrix 9 adding FA to column 20 
	-- signal N10_0_20 : std_logic;
	-- signal N10_1_21 : std_logic;
	FA2517 : full_adder port map (N8_3_20,N9_0_20,N9_1_20,N10_0_20,N10_1_21);
-- In matrix 9 adding FA to column 21 
	-- signal N10_0_21 : std_logic;
	-- signal N10_1_22 : std_logic;
	FA2518 : full_adder port map (N8_3_21,N9_0_21,N9_1_21,N10_0_21,N10_1_22);
-- In matrix 9 adding FA to column 22 
	-- signal N10_0_22 : std_logic;
	-- signal N10_1_23 : std_logic;
	FA2519 : full_adder port map (N8_3_22,N9_0_22,N9_1_22,N10_0_22,N10_1_23);
-- In matrix 9 adding FA to column 23 
	-- signal N10_0_23 : std_logic;
	-- signal N10_1_24 : std_logic;
	FA2520 : full_adder port map (N8_3_23,N9_0_23,N9_1_23,N10_0_23,N10_1_24);
-- In matrix 9 adding FA to column 24 
	-- signal N10_0_24 : std_logic;
	-- signal N10_1_25 : std_logic;
	FA2521 : full_adder port map (N8_3_24,N9_0_24,N9_1_24,N10_0_24,N10_1_25);
-- In matrix 9 adding FA to column 25 
	-- signal N10_0_25 : std_logic;
	-- signal N10_1_26 : std_logic;
	FA2522 : full_adder port map (N8_3_25,N9_0_25,N9_1_25,N10_0_25,N10_1_26);
-- In matrix 9 adding FA to column 26 
	-- signal N10_0_26 : std_logic;
	-- signal N10_1_27 : std_logic;
	FA2523 : full_adder port map (N8_3_26,N9_0_26,N9_1_26,N10_0_26,N10_1_27);
-- In matrix 9 adding FA to column 27 
	-- signal N10_0_27 : std_logic;
	-- signal N10_1_28 : std_logic;
	FA2524 : full_adder port map (N8_3_27,N9_0_27,N9_1_27,N10_0_27,N10_1_28);
-- In matrix 9 adding FA to column 28 
	-- signal N10_0_28 : std_logic;
	-- signal N10_1_29 : std_logic;
	FA2525 : full_adder port map (N8_3_28,N9_0_28,N9_1_28,N10_0_28,N10_1_29);
-- In matrix 9 adding FA to column 29 
	-- signal N10_0_29 : std_logic;
	-- signal N10_1_30 : std_logic;
	FA2526 : full_adder port map (N8_3_29,N9_0_29,N9_1_29,N10_0_29,N10_1_30);
-- In matrix 9 adding FA to column 30 
	-- signal N10_0_30 : std_logic;
	-- signal N10_1_31 : std_logic;
	FA2527 : full_adder port map (N8_3_30,N9_0_30,N9_1_30,N10_0_30,N10_1_31);
-- In matrix 9 adding FA to column 31 
	-- signal N10_0_31 : std_logic;
	-- signal N10_1_32 : std_logic;
	FA2528 : full_adder port map (N8_3_31,N9_0_31,N9_1_31,N10_0_31,N10_1_32);
-- In matrix 9 adding FA to column 32 
	-- signal N10_0_32 : std_logic;
	-- signal N10_1_33 : std_logic;
	FA2529 : full_adder port map (N8_3_32,N9_0_32,N9_1_32,N10_0_32,N10_1_33);
-- In matrix 9 adding FA to column 33 
	-- signal N10_0_33 : std_logic;
	-- signal N10_1_34 : std_logic;
	FA2530 : full_adder port map (N8_3_33,N9_0_33,N9_1_33,N10_0_33,N10_1_34);
-- In matrix 9 adding FA to column 34 
	-- signal N10_0_34 : std_logic;
	-- signal N10_1_35 : std_logic;
	FA2531 : full_adder port map (N8_3_34,N9_0_34,N9_1_34,N10_0_34,N10_1_35);
-- In matrix 9 adding FA to column 35 
	-- signal N10_0_35 : std_logic;
	-- signal N10_1_36 : std_logic;
	FA2532 : full_adder port map (N8_3_35,N9_0_35,N9_1_35,N10_0_35,N10_1_36);
-- In matrix 9 adding FA to column 36 
	-- signal N10_0_36 : std_logic;
	-- signal N10_1_37 : std_logic;
	FA2533 : full_adder port map (N8_3_36,N9_0_36,N9_1_36,N10_0_36,N10_1_37);
-- In matrix 9 adding FA to column 37 
	-- signal N10_0_37 : std_logic;
	-- signal N10_1_38 : std_logic;
	FA2534 : full_adder port map (N8_3_37,N9_0_37,N9_1_37,N10_0_37,N10_1_38);
-- In matrix 9 adding FA to column 38 
	-- signal N10_0_38 : std_logic;
	-- signal N10_1_39 : std_logic;
	FA2535 : full_adder port map (N8_3_38,N9_0_38,N9_1_38,N10_0_38,N10_1_39);
-- In matrix 9 adding FA to column 39 
	-- signal N10_0_39 : std_logic;
	-- signal N10_1_40 : std_logic;
	FA2536 : full_adder port map (N8_3_39,N9_0_39,N9_1_39,N10_0_39,N10_1_40);
-- In matrix 9 adding FA to column 40 
	-- signal N10_0_40 : std_logic;
	-- signal N10_1_41 : std_logic;
	FA2537 : full_adder port map (N8_3_40,N9_0_40,N9_1_40,N10_0_40,N10_1_41);
-- In matrix 9 adding FA to column 41 
	-- signal N10_0_41 : std_logic;
	-- signal N10_1_42 : std_logic;
	FA2538 : full_adder port map (N8_3_41,N9_0_41,N9_1_41,N10_0_41,N10_1_42);
-- In matrix 9 adding FA to column 42 
	-- signal N10_0_42 : std_logic;
	-- signal N10_1_43 : std_logic;
	FA2539 : full_adder port map (N8_3_42,N9_0_42,N9_1_42,N10_0_42,N10_1_43);
-- In matrix 9 adding FA to column 43 
	-- signal N10_0_43 : std_logic;
	-- signal N10_1_44 : std_logic;
	FA2540 : full_adder port map (N8_3_43,N9_0_43,N9_1_43,N10_0_43,N10_1_44);
-- In matrix 9 adding FA to column 44 
	-- signal N10_0_44 : std_logic;
	-- signal N10_1_45 : std_logic;
	FA2541 : full_adder port map (N8_3_44,N9_0_44,N9_1_44,N10_0_44,N10_1_45);
-- In matrix 9 adding FA to column 45 
	-- signal N10_0_45 : std_logic;
	-- signal N10_1_46 : std_logic;
	FA2542 : full_adder port map (N8_3_45,N9_0_45,N9_1_45,N10_0_45,N10_1_46);
-- In matrix 9 adding FA to column 46 
	-- signal N10_0_46 : std_logic;
	-- signal N10_1_47 : std_logic;
	FA2543 : full_adder port map (N8_3_46,N9_0_46,N9_1_46,N10_0_46,N10_1_47);
-- In matrix 9 adding FA to column 47 
	-- signal N10_0_47 : std_logic;
	-- signal N10_1_48 : std_logic;
	FA2544 : full_adder port map (N8_3_47,N9_0_47,N9_1_47,N10_0_47,N10_1_48);
-- In matrix 9 adding FA to column 48 
	-- signal N10_0_48 : std_logic;
	-- signal N10_1_49 : std_logic;
	FA2545 : full_adder port map (N8_3_48,N9_0_48,N9_1_48,N10_0_48,N10_1_49);
-- In matrix 9 adding FA to column 49 
	-- signal N10_0_49 : std_logic;
	-- signal N10_1_50 : std_logic;
	FA2546 : full_adder port map (N8_3_49,N9_0_49,N9_1_49,N10_0_49,N10_1_50);
-- In matrix 9 adding FA to column 50 
	-- signal N10_0_50 : std_logic;
	-- signal N10_1_51 : std_logic;
	FA2547 : full_adder port map (N8_3_50,N9_0_50,N9_1_50,N10_0_50,N10_1_51);
-- In matrix 9 adding FA to column 51 
	-- signal N10_0_51 : std_logic;
	-- signal N10_1_52 : std_logic;
	FA2548 : full_adder port map (N8_3_51,N9_0_51,N9_1_51,N10_0_51,N10_1_52);
-- In matrix 9 adding FA to column 52 
	-- signal N10_0_52 : std_logic;
	-- signal N10_1_53 : std_logic;
	FA2549 : full_adder port map (N8_3_52,N9_0_52,N9_1_52,N10_0_52,N10_1_53);
-- In matrix 9 adding FA to column 53 
	-- signal N10_0_53 : std_logic;
	-- signal N10_1_54 : std_logic;
	FA2550 : full_adder port map (N8_3_53,N9_0_53,N9_1_53,N10_0_53,N10_1_54);
-- In matrix 9 adding FA to column 54 
	-- signal N10_0_54 : std_logic;
	-- signal N10_1_55 : std_logic;
	FA2551 : full_adder port map (N8_3_54,N9_0_54,N9_1_54,N10_0_54,N10_1_55);
-- In matrix 9 adding FA to column 55 
	-- signal N10_0_55 : std_logic;
	-- signal N10_1_56 : std_logic;
	FA2552 : full_adder port map (N8_3_55,N9_0_55,N9_1_55,N10_0_55,N10_1_56);
-- In matrix 9 adding FA to column 56 
	-- signal N10_0_56 : std_logic;
	-- signal N10_1_57 : std_logic;
	FA2553 : full_adder port map (N8_3_56,N9_0_56,N9_1_56,N10_0_56,N10_1_57);
-- In matrix 9 adding FA to column 57 
	-- signal N10_0_57 : std_logic;
	-- signal N10_1_58 : std_logic;
	FA2554 : full_adder port map (N8_3_57,N9_0_57,N9_1_57,N10_0_57,N10_1_58);
-- In matrix 9 adding FA to column 58 
	-- signal N10_0_58 : std_logic;
	-- signal N10_1_59 : std_logic;
	FA2555 : full_adder port map (N8_3_58,N9_0_58,N9_1_58,N10_0_58,N10_1_59);
-- In matrix 9 adding FA to column 59 
	-- signal N10_0_59 : std_logic;
	-- signal N10_1_60 : std_logic;
	FA2556 : full_adder port map (N8_3_59,N9_0_59,N9_1_59,N10_0_59,N10_1_60);
-- In matrix 9 adding FA to column 60 
	-- signal N10_0_60 : std_logic;
	-- signal N10_1_61 : std_logic;
	FA2557 : full_adder port map (N8_3_60,N9_0_60,N9_1_60,N10_0_60,N10_1_61);
-- In matrix 9 adding FA to column 61 
	-- signal N10_0_61 : std_logic;
	-- signal N10_1_62 : std_logic;
	FA2558 : full_adder port map (N8_3_61,N9_0_61,N9_1_61,N10_0_61,N10_1_62);
-- In matrix 9 adding FA to column 62 
	-- signal N10_0_62 : std_logic;
	-- signal N10_1_63 : std_logic;
	FA2559 : full_adder port map (N8_3_62,N9_0_62,N9_1_62,N10_0_62,N10_1_63);
-- In matrix 9 adding FA to column 63 
	-- signal N10_0_63 : std_logic;
	-- signal N10_1_64 : std_logic;
	FA2560 : full_adder port map (N8_3_63,N9_0_63,N9_1_63,N10_0_63,N10_1_64);
-- In matrix 9 adding FA to column 64 
	-- signal N10_0_64 : std_logic;
	-- signal N10_1_65 : std_logic;
	FA2561 : full_adder port map (N8_3_64,N9_0_64,N9_1_64,N10_0_64,N10_1_65);
-- In matrix 9 adding FA to column 65 
	-- signal N10_0_65 : std_logic;
	-- signal N10_1_66 : std_logic;
	FA2562 : full_adder port map (N8_3_65,N9_0_65,N9_1_65,N10_0_65,N10_1_66);
-- In matrix 9 adding FA to column 66 
	-- signal N10_0_66 : std_logic;
	-- signal N10_1_67 : std_logic;
	FA2563 : full_adder port map (N8_3_66,N9_0_66,N9_1_66,N10_0_66,N10_1_67);
-- In matrix 9 adding FA to column 67 
	-- signal N10_0_67 : std_logic;
	-- signal N10_1_68 : std_logic;
	FA2564 : full_adder port map (N8_3_67,N9_0_67,N9_1_67,N10_0_67,N10_1_68);
-- In matrix 9 adding FA to column 68 
	-- signal N10_0_68 : std_logic;
	-- signal N10_1_69 : std_logic;
	FA2565 : full_adder port map (N8_3_68,N9_0_68,N9_1_68,N10_0_68,N10_1_69);
-- In matrix 9 adding FA to column 69 
	-- signal N10_0_69 : std_logic;
	-- signal N10_1_70 : std_logic;
	FA2566 : full_adder port map (N8_3_69,N9_0_69,N9_1_69,N10_0_69,N10_1_70);
-- In matrix 9 adding FA to column 70 
	-- signal N10_0_70 : std_logic;
	-- signal N10_1_71 : std_logic;
	FA2567 : full_adder port map (N8_3_70,N9_0_70,N9_1_70,N10_0_70,N10_1_71);
-- In matrix 9 adding FA to column 71 
	-- signal N10_0_71 : std_logic;
	-- signal N10_1_72 : std_logic;
	FA2568 : full_adder port map (N8_3_71,N9_0_71,N9_1_71,N10_0_71,N10_1_72);
-- In matrix 9 adding FA to column 72 
	-- signal N10_0_72 : std_logic;
	-- signal N10_1_73 : std_logic;
	FA2569 : full_adder port map (N8_3_72,N9_0_72,N9_1_72,N10_0_72,N10_1_73);
-- In matrix 9 adding FA to column 73 
	-- signal N10_0_73 : std_logic;
	-- signal N10_1_74 : std_logic;
	FA2570 : full_adder port map (N8_3_73,N9_0_73,N9_1_73,N10_0_73,N10_1_74);
-- In matrix 9 adding FA to column 74 
	-- signal N10_0_74 : std_logic;
	-- signal N10_1_75 : std_logic;
	FA2571 : full_adder port map (N8_3_74,N9_0_74,N9_1_74,N10_0_74,N10_1_75);
-- In matrix 9 adding FA to column 75 
	-- signal N10_0_75 : std_logic;
	-- signal N10_1_76 : std_logic;
	FA2572 : full_adder port map (N8_3_75,N9_0_75,N9_1_75,N10_0_75,N10_1_76);
-- In matrix 9 adding FA to column 76 
	-- signal N10_0_76 : std_logic;
	-- signal N10_1_77 : std_logic;
	FA2573 : full_adder port map (N8_3_76,N9_0_76,N9_1_76,N10_0_76,N10_1_77);
-- In matrix 9 adding FA to column 77 
	-- signal N10_0_77 : std_logic;
	-- signal N10_1_78 : std_logic;
	FA2574 : full_adder port map (N8_3_77,N9_0_77,N9_1_77,N10_0_77,N10_1_78);
-- In matrix 9 adding FA to column 78 
	-- signal N10_0_78 : std_logic;
	-- signal N10_1_79 : std_logic;
	FA2575 : full_adder port map (N8_3_78,N9_0_78,N9_1_78,N10_0_78,N10_1_79);
-- In matrix 9 adding FA to column 79 
	-- signal N10_0_79 : std_logic;
	-- signal N10_1_80 : std_logic;
	FA2576 : full_adder port map (N8_3_79,N9_0_79,N9_1_79,N10_0_79,N10_1_80);
-- In matrix 9 adding FA to column 80 
	-- signal N10_0_80 : std_logic;
	-- signal N10_1_81 : std_logic;
	FA2577 : full_adder port map (N8_3_80,N9_0_80,N9_1_80,N10_0_80,N10_1_81);
-- In matrix 9 adding FA to column 81 
	-- signal N10_0_81 : std_logic;
	-- signal N10_1_82 : std_logic;
	FA2578 : full_adder port map (N8_3_81,N9_0_81,N9_1_81,N10_0_81,N10_1_82);
-- In matrix 9 adding FA to column 82 
	-- signal N10_0_82 : std_logic;
	-- signal N10_1_83 : std_logic;
	FA2579 : full_adder port map (N8_3_82,N9_0_82,N9_1_82,N10_0_82,N10_1_83);
-- In matrix 9 adding FA to column 83 
	-- signal N10_0_83 : std_logic;
	-- signal N10_1_84 : std_logic;
	FA2580 : full_adder port map (N8_3_83,N9_0_83,N9_1_83,N10_0_83,N10_1_84);
-- In matrix 9 adding FA to column 84 
	-- signal N10_0_84 : std_logic;
	-- signal N10_1_85 : std_logic;
	FA2581 : full_adder port map (N8_3_84,N9_0_84,N9_1_84,N10_0_84,N10_1_85);
-- In matrix 9 adding FA to column 85 
	-- signal N10_0_85 : std_logic;
	-- signal N10_1_86 : std_logic;
	FA2582 : full_adder port map (N8_3_85,N9_0_85,N9_1_85,N10_0_85,N10_1_86);
-- In matrix 9 adding FA to column 86 
	-- signal N10_0_86 : std_logic;
	-- signal N10_1_87 : std_logic;
	FA2583 : full_adder port map (N8_3_86,N9_0_86,N9_1_86,N10_0_86,N10_1_87);
-- In matrix 9 adding FA to column 87 
	-- signal N10_0_87 : std_logic;
	-- signal N10_1_88 : std_logic;
	FA2584 : full_adder port map (N8_3_87,N9_0_87,N9_1_87,N10_0_87,N10_1_88);
-- In matrix 9 adding FA to column 88 
	-- signal N10_0_88 : std_logic;
	-- signal N10_1_89 : std_logic;
	FA2585 : full_adder port map (N8_3_88,N9_0_88,N9_1_88,N10_0_88,N10_1_89);
-- In matrix 9 adding FA to column 89 
	-- signal N10_0_89 : std_logic;
	-- signal N10_1_90 : std_logic;
	FA2586 : full_adder port map (N8_3_89,N9_0_89,N9_1_89,N10_0_89,N10_1_90);
-- In matrix 9 adding FA to column 90 
	-- signal N10_0_90 : std_logic;
	-- signal N10_1_91 : std_logic;
	FA2587 : full_adder port map (N8_3_90,N9_0_90,N9_1_90,N10_0_90,N10_1_91);
-- In matrix 9 adding FA to column 91 
	-- signal N10_0_91 : std_logic;
	-- signal N10_1_92 : std_logic;
	FA2588 : full_adder port map (N8_3_91,N9_0_91,N9_1_91,N10_0_91,N10_1_92);
-- In matrix 9 adding FA to column 92 
	-- signal N10_0_92 : std_logic;
	-- signal N10_1_93 : std_logic;
	FA2589 : full_adder port map (N8_3_92,N9_0_92,N9_1_92,N10_0_92,N10_1_93);
-- In matrix 9 adding FA to column 93 
	-- signal N10_0_93 : std_logic;
	-- signal N10_1_94 : std_logic;
	FA2590 : full_adder port map (N8_3_93,N9_0_93,N9_1_93,N10_0_93,N10_1_94);
-- In matrix 9 adding FA to column 94 
	-- signal N10_0_94 : std_logic;
	-- signal N10_1_95 : std_logic;
	FA2591 : full_adder port map (N8_3_94,N9_0_94,N9_1_94,N10_0_94,N10_1_95);
-- In matrix 9 adding FA to column 95 
	-- signal N10_0_95 : std_logic;
	-- signal N10_1_96 : std_logic;
	FA2592 : full_adder port map (N8_3_95,N9_0_95,N9_1_95,N10_0_95,N10_1_96);
-- In matrix 9 adding FA to column 96 
	-- signal N10_0_96 : std_logic;
	-- signal N10_1_97 : std_logic;
	FA2593 : full_adder port map (N8_3_96,N9_0_96,N9_1_96,N10_0_96,N10_1_97);
-- In matrix 9 adding FA to column 97 
	-- signal N10_0_97 : std_logic;
	-- signal N10_1_98 : std_logic;
	FA2594 : full_adder port map (N8_3_97,N9_0_97,N9_1_97,N10_0_97,N10_1_98);
-- In matrix 9 adding FA to column 98 
	-- signal N10_0_98 : std_logic;
	-- signal N10_1_99 : std_logic;
	FA2595 : full_adder port map (N8_3_98,N9_0_98,N9_1_98,N10_0_98,N10_1_99);
-- In matrix 9 adding FA to column 99 
	-- signal N10_0_99 : std_logic;
	-- signal N10_1_100 : std_logic;
	FA2596 : full_adder port map (N8_3_99,N9_0_99,N9_1_99,N10_0_99,N10_1_100);
-- In matrix 9 adding FA to column 100 
	-- signal N10_0_100 : std_logic;
	-- signal N10_1_101 : std_logic;
	FA2597 : full_adder port map (N8_3_100,N9_0_100,N9_1_100,N10_0_100,N10_1_101);
-- In matrix 9 adding FA to column 101 
	-- signal N10_0_101 : std_logic;
	-- signal N10_1_102 : std_logic;
	FA2598 : full_adder port map (N8_3_101,N9_0_101,N9_1_101,N10_0_101,N10_1_102);
-- In matrix 9 adding FA to column 102 
	-- signal N10_0_102 : std_logic;
	-- signal N10_1_103 : std_logic;
	FA2599 : full_adder port map (N8_1_102,N9_0_102,N9_1_102,N10_0_102,N10_1_103);
-- In matrix 9 adding FA to column 103 
	-- signal N10_0_103 : std_logic;
	-- signal N10_1_104 : std_logic;
	FA2600 : full_adder port map (N0_51_103,N0_52_103,N9_1_103,N10_0_103,N10_1_104);

	S(0) <= '0';
	S(1) <= N0_0_1;
	S(2) <= N0_2_2;
	S(3) <= N10_0_3;
	S(4) <= N10_0_4;
	S(5) <= N10_0_5;
	S(6) <= N10_0_6;
	S(7) <= N10_0_7;
	S(8) <= N10_0_8;
	S(9) <= N10_0_9;
	S(10) <= N10_0_10;
	S(11) <= N10_0_11;
	S(12) <= N10_0_12;
	S(13) <= N10_0_13;
	S(14) <= N10_0_14;
	S(15) <= N10_0_15;
	S(16) <= N10_0_16;
	S(17) <= N10_0_17;
	S(18) <= N10_0_18;
	S(19) <= N10_0_19;
	S(20) <= N10_0_20;
	S(21) <= N10_0_21;
	S(22) <= N10_0_22;
	S(23) <= N10_0_23;
	S(24) <= N10_0_24;
	S(25) <= N10_0_25;
	S(26) <= N10_0_26;
	S(27) <= N10_0_27;
	S(28) <= N10_0_28;
	S(29) <= N10_0_29;
	S(30) <= N10_0_30;
	S(31) <= N10_0_31;
	S(32) <= N10_0_32;
	S(33) <= N10_0_33;
	S(34) <= N10_0_34;
	S(35) <= N10_0_35;
	S(36) <= N10_0_36;
	S(37) <= N10_0_37;
	S(38) <= N10_0_38;
	S(39) <= N10_0_39;
	S(40) <= N10_0_40;
	S(41) <= N10_0_41;
	S(42) <= N10_0_42;
	S(43) <= N10_0_43;
	S(44) <= N10_0_44;
	S(45) <= N10_0_45;
	S(46) <= N10_0_46;
	S(47) <= N10_0_47;
	S(48) <= N10_0_48;
	S(49) <= N10_0_49;
	S(50) <= N10_0_50;
	S(51) <= N10_0_51;
	S(52) <= N10_0_52;
	S(53) <= N10_0_53;
	S(54) <= N10_0_54;
	S(55) <= N10_0_55;
	S(56) <= N10_0_56;
	S(57) <= N10_0_57;
	S(58) <= N10_0_58;
	S(59) <= N10_0_59;
	S(60) <= N10_0_60;
	S(61) <= N10_0_61;
	S(62) <= N10_0_62;
	S(63) <= N10_0_63;
	S(64) <= N10_0_64;
	S(65) <= N10_0_65;
	S(66) <= N10_0_66;
	S(67) <= N10_0_67;
	S(68) <= N10_0_68;
	S(69) <= N10_0_69;
	S(70) <= N10_0_70;
	S(71) <= N10_0_71;
	S(72) <= N10_0_72;
	S(73) <= N10_0_73;
	S(74) <= N10_0_74;
	S(75) <= N10_0_75;
	S(76) <= N10_0_76;
	S(77) <= N10_0_77;
	S(78) <= N10_0_78;
	S(79) <= N10_0_79;
	S(80) <= N10_0_80;
	S(81) <= N10_0_81;
	S(82) <= N10_0_82;
	S(83) <= N10_0_83;
	S(84) <= N10_0_84;
	S(85) <= N10_0_85;
	S(86) <= N10_0_86;
	S(87) <= N10_0_87;
	S(88) <= N10_0_88;
	S(89) <= N10_0_89;
	S(90) <= N10_0_90;
	S(91) <= N10_0_91;
	S(92) <= N10_0_92;
	S(93) <= N10_0_93;
	S(94) <= N10_0_94;
	S(95) <= N10_0_95;
	S(96) <= N10_0_96;
	S(97) <= N10_0_97;
	S(98) <= N10_0_98;
	S(99) <= N10_0_99;
	S(100) <= N10_0_100;
	S(101) <= N10_0_101;
	S(102) <= N10_0_102;
	S(103) <= N10_0_103;
	S(104) <= N0_52_104;
        S(105) <= '0';
        
	C(0) <= N0_0_0;
	C(1) <= N0_1_1;
	C(2) <= N10_0_2;
	C(3) <= N10_1_3;
	C(4) <= N10_1_4;
	C(5) <= N10_1_5;
	C(6) <= N10_1_6;
	C(7) <= N10_1_7;
	C(8) <= N10_1_8;
	C(9) <= N10_1_9;
	C(10) <= N10_1_10;
	C(11) <= N10_1_11;
	C(12) <= N10_1_12;
	C(13) <= N10_1_13;
	C(14) <= N10_1_14;
	C(15) <= N10_1_15;
	C(16) <= N10_1_16;
	C(17) <= N10_1_17;
	C(18) <= N10_1_18;
	C(19) <= N10_1_19;
	C(20) <= N10_1_20;
	C(21) <= N10_1_21;
	C(22) <= N10_1_22;
	C(23) <= N10_1_23;
	C(24) <= N10_1_24;
	C(25) <= N10_1_25;
	C(26) <= N10_1_26;
	C(27) <= N10_1_27;
	C(28) <= N10_1_28;
	C(29) <= N10_1_29;
	C(30) <= N10_1_30;
	C(31) <= N10_1_31;
	C(32) <= N10_1_32;
	C(33) <= N10_1_33;
	C(34) <= N10_1_34;
	C(35) <= N10_1_35;
	C(36) <= N10_1_36;
	C(37) <= N10_1_37;
	C(38) <= N10_1_38;
	C(39) <= N10_1_39;
	C(40) <= N10_1_40;
	C(41) <= N10_1_41;
	C(42) <= N10_1_42;
	C(43) <= N10_1_43;
	C(44) <= N10_1_44;
	C(45) <= N10_1_45;
	C(46) <= N10_1_46;
	C(47) <= N10_1_47;
	C(48) <= N10_1_48;
	C(49) <= N10_1_49;
	C(50) <= N10_1_50;
	C(51) <= N10_1_51;
	C(52) <= N10_1_52;
	C(53) <= N10_1_53;
	C(54) <= N10_1_54;
	C(55) <= N10_1_55;
	C(56) <= N10_1_56;
	C(57) <= N10_1_57;
	C(58) <= N10_1_58;
	C(59) <= N10_1_59;
	C(60) <= N10_1_60;
	C(61) <= N10_1_61;
	C(62) <= N10_1_62;
	C(63) <= N10_1_63;
	C(64) <= N10_1_64;
	C(65) <= N10_1_65;
	C(66) <= N10_1_66;
	C(67) <= N10_1_67;
	C(68) <= N10_1_68;
	C(69) <= N10_1_69;
	C(70) <= N10_1_70;
	C(71) <= N10_1_71;
	C(72) <= N10_1_72;
	C(73) <= N10_1_73;
	C(74) <= N10_1_74;
	C(75) <= N10_1_75;
	C(76) <= N10_1_76;
	C(77) <= N10_1_77;
	C(78) <= N10_1_78;
	C(79) <= N10_1_79;
	C(80) <= N10_1_80;
	C(81) <= N10_1_81;
	C(82) <= N10_1_82;
	C(83) <= N10_1_83;
	C(84) <= N10_1_84;
	C(85) <= N10_1_85;
	C(86) <= N10_1_86;
	C(87) <= N10_1_87;
	C(88) <= N10_1_88;
	C(89) <= N10_1_89;
	C(90) <= N10_1_90;
	C(91) <= N10_1_91;
	C(92) <= N10_1_92;
	C(93) <= N10_1_93;
	C(94) <= N10_1_94;
	C(95) <= N10_1_95;
	C(96) <= N10_1_96;
	C(97) <= N10_1_97;
	C(98) <= N10_1_98;
	C(99) <= N10_1_99;
	C(100) <= N10_1_100;
	C(101) <= N10_1_101;
	C(102) <= N10_1_102;
	C(103) <= N10_1_103;
	C(104) <= N10_1_104;
        C(105) <= '0';
        
end Structure;

